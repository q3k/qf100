magic
tech sky130A
magscale 1 2
timestamp 1647787628
<< viali >>
rect 1593 47209 1627 47243
rect 3065 47209 3099 47243
rect 5457 47209 5491 47243
rect 6561 47209 6595 47243
rect 7297 47209 7331 47243
rect 8125 47209 8159 47243
rect 9137 47209 9171 47243
rect 9873 47209 9907 47243
rect 10609 47209 10643 47243
rect 11713 47209 11747 47243
rect 12449 47209 12483 47243
rect 13185 47209 13219 47243
rect 14289 47209 14323 47243
rect 15025 47209 15059 47243
rect 15761 47209 15795 47243
rect 17601 47209 17635 47243
rect 18337 47209 18371 47243
rect 20177 47209 20211 47243
rect 20913 47209 20947 47243
rect 22293 47209 22327 47243
rect 23121 47209 23155 47243
rect 24593 47209 24627 47243
rect 26065 47209 26099 47243
rect 27537 47209 27571 47243
rect 35357 47209 35391 47243
rect 4721 47141 4755 47175
rect 31309 47141 31343 47175
rect 28365 47073 28399 47107
rect 29561 47073 29595 47107
rect 35909 47073 35943 47107
rect 37289 47073 37323 47107
rect 1409 47005 1443 47039
rect 2145 47005 2179 47039
rect 2881 47005 2915 47039
rect 3801 47005 3835 47039
rect 4537 47005 4571 47039
rect 5273 47005 5307 47039
rect 6377 47005 6411 47039
rect 7113 47005 7147 47039
rect 7941 47005 7975 47039
rect 8953 47005 8987 47039
rect 9689 47005 9723 47039
rect 10425 47005 10459 47039
rect 11529 47005 11563 47039
rect 12265 47005 12299 47039
rect 13001 47005 13035 47039
rect 14105 47005 14139 47039
rect 14841 47005 14875 47039
rect 15577 47005 15611 47039
rect 16681 47005 16715 47039
rect 17417 47005 17451 47039
rect 18153 47005 18187 47039
rect 19257 47005 19291 47039
rect 19993 47005 20027 47039
rect 20729 47005 20763 47039
rect 22109 47005 22143 47039
rect 22937 47005 22971 47039
rect 24409 47005 24443 47039
rect 25145 47005 25179 47039
rect 25881 47005 25915 47039
rect 27445 47005 27479 47039
rect 29837 47005 29871 47039
rect 31493 47005 31527 47039
rect 32137 47005 32171 47039
rect 32413 47005 32447 47039
rect 33885 47005 33919 47039
rect 35265 47005 35299 47039
rect 36185 47005 36219 47039
rect 37565 47005 37599 47039
rect 28181 46937 28215 46971
rect 34069 46937 34103 46971
rect 2329 46869 2363 46903
rect 3985 46869 4019 46903
rect 16865 46869 16899 46903
rect 19441 46869 19475 46903
rect 25329 46869 25363 46903
rect 5641 46665 5675 46699
rect 12173 46665 12207 46699
rect 14289 46665 14323 46699
rect 15945 46665 15979 46699
rect 17693 46665 17727 46699
rect 18521 46665 18555 46699
rect 19533 46665 19567 46699
rect 21005 46665 21039 46699
rect 23857 46665 23891 46699
rect 27169 46665 27203 46699
rect 13829 46597 13863 46631
rect 17049 46597 17083 46631
rect 34713 46597 34747 46631
rect 5457 46529 5491 46563
rect 12357 46529 12391 46563
rect 13001 46529 13035 46563
rect 13645 46529 13679 46563
rect 14473 46529 14507 46563
rect 15485 46529 15519 46563
rect 16129 46529 16163 46563
rect 16865 46529 16899 46563
rect 17325 46529 17359 46563
rect 17877 46529 17911 46563
rect 18705 46529 18739 46563
rect 19717 46529 19751 46563
rect 21189 46529 21223 46563
rect 21833 46529 21867 46563
rect 24041 46529 24075 46563
rect 26985 46529 27019 46563
rect 29653 46529 29687 46563
rect 32321 46529 32355 46563
rect 33149 46529 33183 46563
rect 37289 46529 37323 46563
rect 13461 46461 13495 46495
rect 16681 46461 16715 46495
rect 29929 46461 29963 46495
rect 37565 46461 37599 46495
rect 12817 46393 12851 46427
rect 15301 46393 15335 46427
rect 22017 46393 22051 46427
rect 32137 46325 32171 46359
rect 32965 46325 32999 46359
rect 34805 46325 34839 46359
rect 12265 46121 12299 46155
rect 13461 46121 13495 46155
rect 14841 46121 14875 46155
rect 16497 46121 16531 46155
rect 17785 46121 17819 46155
rect 22201 46121 22235 46155
rect 15669 46053 15703 46087
rect 13093 45985 13127 46019
rect 16129 45985 16163 46019
rect 11989 45917 12023 45951
rect 12081 45917 12115 45951
rect 13277 45917 13311 45951
rect 14473 45917 14507 45951
rect 14657 45917 14691 45951
rect 15301 45917 15335 45951
rect 15485 45917 15519 45951
rect 16313 45917 16347 45951
rect 17049 45917 17083 45951
rect 17141 45917 17175 45951
rect 17325 45917 17359 45951
rect 17969 45917 18003 45951
rect 22385 45917 22419 45951
rect 37197 45917 37231 45951
rect 37933 45917 37967 45951
rect 37289 45781 37323 45815
rect 38025 45781 38059 45815
rect 23305 45577 23339 45611
rect 17693 45509 17727 45543
rect 20177 45509 20211 45543
rect 21281 45509 21315 45543
rect 22661 45509 22695 45543
rect 13093 45441 13127 45475
rect 13829 45441 13863 45475
rect 17509 45441 17543 45475
rect 19349 45441 19383 45475
rect 19993 45441 20027 45475
rect 21097 45441 21131 45475
rect 22477 45441 22511 45475
rect 23213 45441 23247 45475
rect 29745 45441 29779 45475
rect 13553 45373 13587 45407
rect 17325 45373 17359 45407
rect 19809 45373 19843 45407
rect 20913 45373 20947 45407
rect 22293 45373 22327 45407
rect 12909 45305 12943 45339
rect 19165 45305 19199 45339
rect 29929 45305 29963 45339
rect 22937 45237 22971 45271
rect 21373 45033 21407 45067
rect 17877 44897 17911 44931
rect 19625 44897 19659 44931
rect 23305 44897 23339 44931
rect 18153 44829 18187 44863
rect 19349 44829 19383 44863
rect 23029 44829 23063 44863
rect 21281 44761 21315 44795
rect 16129 44489 16163 44523
rect 18337 44489 18371 44523
rect 23857 44489 23891 44523
rect 13176 44353 13210 44387
rect 15005 44353 15039 44387
rect 18153 44353 18187 44387
rect 20076 44353 20110 44387
rect 22845 44353 22879 44387
rect 24041 44353 24075 44387
rect 12909 44285 12943 44319
rect 14749 44285 14783 44319
rect 17969 44285 18003 44319
rect 19809 44285 19843 44319
rect 22569 44285 22603 44319
rect 14289 44149 14323 44183
rect 21189 44149 21223 44183
rect 20637 43945 20671 43979
rect 23305 43945 23339 43979
rect 17785 43809 17819 43843
rect 14289 43741 14323 43775
rect 15669 43741 15703 43775
rect 17509 43741 17543 43775
rect 19257 43741 19291 43775
rect 20913 43741 20947 43775
rect 22937 43741 22971 43775
rect 23121 43741 23155 43775
rect 14105 43673 14139 43707
rect 15914 43673 15948 43707
rect 19502 43673 19536 43707
rect 21158 43673 21192 43707
rect 22661 43673 22695 43707
rect 14473 43605 14507 43639
rect 17049 43605 17083 43639
rect 22293 43605 22327 43639
rect 14105 43401 14139 43435
rect 14565 43401 14599 43435
rect 23949 43401 23983 43435
rect 24593 43401 24627 43435
rect 20085 43333 20119 43367
rect 12725 43265 12759 43299
rect 12992 43265 13026 43299
rect 14795 43265 14829 43299
rect 14933 43265 14967 43299
rect 15025 43265 15059 43299
rect 15209 43265 15243 43299
rect 15761 43265 15795 43299
rect 15945 43265 15979 43299
rect 16681 43265 16715 43299
rect 16937 43265 16971 43299
rect 19901 43265 19935 43299
rect 24133 43265 24167 43299
rect 24777 43265 24811 43299
rect 16129 43061 16163 43095
rect 18061 43061 18095 43095
rect 20269 43061 20303 43095
rect 15577 42857 15611 42891
rect 24777 42857 24811 42891
rect 20545 42789 20579 42823
rect 14105 42721 14139 42755
rect 22017 42721 22051 42755
rect 25053 42721 25087 42755
rect 13369 42653 13403 42687
rect 14381 42653 14415 42687
rect 14473 42653 14507 42687
rect 14565 42653 14599 42687
rect 14749 42653 14783 42687
rect 15853 42653 15887 42687
rect 15945 42653 15979 42687
rect 16037 42653 16071 42687
rect 16221 42653 16255 42687
rect 19533 42653 19567 42687
rect 20821 42653 20855 42687
rect 20910 42653 20944 42687
rect 21026 42653 21060 42687
rect 21189 42653 21223 42687
rect 24409 42653 24443 42687
rect 24593 42653 24627 42687
rect 13185 42585 13219 42619
rect 13553 42585 13587 42619
rect 19349 42585 19383 42619
rect 21649 42585 21683 42619
rect 21833 42585 21867 42619
rect 22477 42585 22511 42619
rect 22661 42585 22695 42619
rect 19717 42517 19751 42551
rect 22845 42517 22879 42551
rect 14197 42313 14231 42347
rect 15301 42313 15335 42347
rect 17509 42313 17543 42347
rect 19073 42313 19107 42347
rect 20177 42313 20211 42347
rect 24225 42313 24259 42347
rect 14427 42177 14461 42211
rect 14578 42177 14612 42211
rect 14678 42177 14712 42211
rect 14841 42177 14875 42211
rect 15531 42177 15565 42211
rect 15666 42177 15700 42211
rect 15761 42177 15795 42211
rect 15945 42177 15979 42211
rect 18153 42177 18187 42211
rect 19303 42177 19337 42211
rect 19441 42177 19475 42211
rect 19533 42177 19567 42211
rect 19717 42177 19751 42211
rect 20453 42177 20487 42211
rect 20545 42177 20579 42211
rect 20637 42177 20671 42211
rect 20821 42177 20855 42211
rect 22017 42177 22051 42211
rect 22273 42177 22307 42211
rect 24041 42177 24075 42211
rect 17049 42109 17083 42143
rect 23857 42109 23891 42143
rect 17325 42041 17359 42075
rect 17969 41973 18003 42007
rect 23397 41973 23431 42007
rect 17141 41769 17175 41803
rect 22569 41769 22603 41803
rect 27537 41769 27571 41803
rect 14381 41633 14415 41667
rect 13553 41565 13587 41599
rect 14105 41565 14139 41599
rect 19625 41565 19659 41599
rect 19901 41565 19935 41599
rect 15853 41497 15887 41531
rect 21281 41497 21315 41531
rect 27445 41497 27479 41531
rect 13369 41429 13403 41463
rect 15117 41225 15151 41259
rect 15485 41225 15519 41259
rect 17233 41225 17267 41259
rect 12725 41157 12759 41191
rect 12941 41157 12975 41191
rect 14749 41157 14783 41191
rect 15761 41157 15795 41191
rect 15977 41157 16011 41191
rect 17049 41157 17083 41191
rect 17960 41157 17994 41191
rect 22170 41157 22204 41191
rect 14933 41089 14967 41123
rect 17693 41089 17727 41123
rect 13553 41021 13587 41055
rect 13829 41021 13863 41055
rect 19533 41021 19567 41055
rect 19809 41021 19843 41055
rect 21925 41021 21959 41055
rect 12449 40953 12483 40987
rect 16681 40953 16715 40987
rect 23305 40953 23339 40987
rect 12909 40885 12943 40919
rect 13093 40885 13127 40919
rect 15945 40885 15979 40919
rect 16129 40885 16163 40919
rect 17049 40885 17083 40919
rect 19073 40885 19107 40919
rect 12265 40681 12299 40715
rect 13093 40681 13127 40715
rect 16865 40681 16899 40715
rect 18061 40681 18095 40715
rect 20637 40681 20671 40715
rect 12173 40613 12207 40647
rect 14657 40545 14691 40579
rect 12725 40477 12759 40511
rect 16497 40477 16531 40511
rect 16681 40477 16715 40511
rect 17325 40477 17359 40511
rect 17509 40477 17543 40511
rect 17969 40477 18003 40511
rect 18153 40477 18187 40511
rect 19625 40477 19659 40511
rect 20867 40477 20901 40511
rect 21002 40477 21036 40511
rect 21097 40477 21131 40511
rect 21281 40477 21315 40511
rect 22109 40477 22143 40511
rect 22201 40477 22235 40511
rect 22298 40477 22332 40511
rect 22477 40477 22511 40511
rect 11805 40409 11839 40443
rect 14924 40409 14958 40443
rect 17417 40409 17451 40443
rect 21833 40409 21867 40443
rect 13093 40341 13127 40375
rect 13277 40341 13311 40375
rect 16037 40341 16071 40375
rect 19441 40341 19475 40375
rect 19257 40137 19291 40171
rect 24149 40137 24183 40171
rect 15485 40069 15519 40103
rect 15669 40069 15703 40103
rect 19901 40069 19935 40103
rect 20101 40069 20135 40103
rect 20913 40069 20947 40103
rect 21097 40069 21131 40103
rect 23949 40069 23983 40103
rect 11805 40001 11839 40035
rect 12817 40001 12851 40035
rect 13084 40001 13118 40035
rect 14841 40001 14875 40035
rect 18337 40001 18371 40035
rect 18521 40001 18555 40035
rect 18797 40001 18831 40035
rect 21281 40001 21315 40035
rect 24869 40001 24903 40035
rect 25053 40001 25087 40035
rect 11529 39933 11563 39967
rect 18429 39933 18463 39967
rect 23029 39933 23063 39967
rect 14657 39865 14691 39899
rect 19165 39865 19199 39899
rect 19625 39865 19659 39899
rect 23305 39865 23339 39899
rect 23489 39865 23523 39899
rect 14197 39797 14231 39831
rect 15853 39797 15887 39831
rect 20085 39797 20119 39831
rect 20269 39797 20303 39831
rect 24133 39797 24167 39831
rect 24317 39797 24351 39831
rect 12541 39593 12575 39627
rect 13277 39593 13311 39627
rect 14933 39593 14967 39627
rect 25237 39593 25271 39627
rect 25513 39593 25547 39627
rect 26065 39593 26099 39627
rect 25145 39525 25179 39559
rect 16037 39457 16071 39491
rect 11621 39389 11655 39423
rect 12541 39389 12575 39423
rect 12725 39389 12759 39423
rect 13185 39389 13219 39423
rect 13369 39389 13403 39423
rect 15209 39389 15243 39423
rect 15301 39389 15335 39423
rect 15393 39389 15427 39423
rect 15577 39389 15611 39423
rect 19441 39389 19475 39423
rect 19901 39389 19935 39423
rect 21925 39389 21959 39423
rect 16282 39321 16316 39355
rect 17877 39321 17911 39355
rect 18061 39321 18095 39355
rect 21005 39321 21039 39355
rect 21189 39321 21223 39355
rect 22192 39321 22226 39355
rect 24777 39321 24811 39355
rect 25881 39321 25915 39355
rect 11437 39253 11471 39287
rect 17417 39253 17451 39287
rect 18245 39253 18279 39287
rect 19257 39253 19291 39287
rect 20545 39253 20579 39287
rect 21373 39253 21407 39287
rect 23305 39253 23339 39287
rect 26081 39253 26115 39287
rect 26249 39253 26283 39287
rect 12081 39049 12115 39083
rect 15485 39049 15519 39083
rect 21189 39049 21223 39083
rect 26249 39049 26283 39083
rect 22630 38981 22664 39015
rect 24676 38981 24710 39015
rect 15761 38913 15795 38947
rect 15853 38913 15887 38947
rect 15945 38913 15979 38947
rect 16129 38913 16163 38947
rect 17509 38913 17543 38947
rect 17765 38913 17799 38947
rect 19809 38913 19843 38947
rect 20076 38913 20110 38947
rect 22385 38913 22419 38947
rect 26433 38913 26467 38947
rect 11621 38845 11655 38879
rect 24409 38845 24443 38879
rect 11897 38777 11931 38811
rect 18889 38709 18923 38743
rect 23765 38709 23799 38743
rect 25789 38709 25823 38743
rect 12725 38505 12759 38539
rect 13277 38505 13311 38539
rect 15853 38505 15887 38539
rect 17325 38505 17359 38539
rect 19809 38505 19843 38539
rect 22109 38505 22143 38539
rect 23213 38505 23247 38539
rect 25513 38505 25547 38539
rect 19993 38437 20027 38471
rect 21005 38437 21039 38471
rect 25145 38437 25179 38471
rect 25697 38437 25731 38471
rect 12357 38369 12391 38403
rect 10701 38301 10735 38335
rect 14289 38301 14323 38335
rect 15669 38301 15703 38335
rect 16313 38301 16347 38335
rect 16589 38301 16623 38335
rect 16681 38301 16715 38335
rect 17601 38301 17635 38335
rect 17693 38301 17727 38335
rect 17785 38301 17819 38335
rect 17969 38301 18003 38335
rect 19441 38301 19475 38335
rect 21281 38301 21315 38335
rect 21373 38301 21407 38335
rect 21465 38301 21499 38335
rect 21649 38301 21683 38335
rect 22385 38301 22419 38335
rect 22477 38301 22511 38335
rect 22569 38301 22603 38335
rect 22753 38301 22787 38335
rect 23213 38301 23247 38335
rect 23397 38301 23431 38335
rect 26157 38301 26191 38335
rect 26341 38301 26375 38335
rect 13093 38233 13127 38267
rect 15485 38233 15519 38267
rect 16497 38233 16531 38267
rect 19809 38233 19843 38267
rect 25513 38233 25547 38267
rect 26249 38233 26283 38267
rect 13293 38165 13327 38199
rect 13461 38165 13495 38199
rect 14105 38165 14139 38199
rect 16865 38165 16899 38199
rect 10701 37961 10735 37995
rect 12909 37961 12943 37995
rect 14289 37961 14323 37995
rect 19441 37961 19475 37995
rect 20085 37961 20119 37995
rect 21189 37961 21223 37995
rect 22201 37961 22235 37995
rect 25237 37961 25271 37995
rect 27721 37961 27755 37995
rect 29393 37961 29427 37995
rect 14105 37893 14139 37927
rect 14749 37893 14783 37927
rect 14949 37893 14983 37927
rect 18521 37893 18555 37927
rect 21833 37893 21867 37927
rect 29193 37893 29227 37927
rect 9321 37825 9355 37859
rect 9588 37825 9622 37859
rect 11529 37825 11563 37859
rect 11785 37825 11819 37859
rect 16681 37825 16715 37859
rect 18245 37825 18279 37859
rect 18429 37825 18463 37859
rect 18613 37825 18647 37859
rect 19349 37825 19383 37859
rect 19533 37825 19567 37859
rect 19993 37825 20027 37859
rect 20177 37825 20211 37859
rect 21097 37825 21131 37859
rect 22017 37825 22051 37859
rect 25145 37825 25179 37859
rect 25329 37825 25363 37859
rect 27629 37825 27663 37859
rect 16957 37757 16991 37791
rect 28273 37757 28307 37791
rect 28733 37757 28767 37791
rect 13737 37689 13771 37723
rect 15117 37689 15151 37723
rect 28549 37689 28583 37723
rect 14105 37621 14139 37655
rect 14933 37621 14967 37655
rect 18797 37621 18831 37655
rect 29377 37621 29411 37655
rect 29561 37621 29595 37655
rect 12081 37417 12115 37451
rect 23673 37417 23707 37451
rect 11713 37349 11747 37383
rect 13369 37349 13403 37383
rect 23305 37349 23339 37383
rect 24961 37349 24995 37383
rect 8953 37281 8987 37315
rect 16037 37281 16071 37315
rect 17693 37281 17727 37315
rect 28917 37281 28951 37315
rect 14105 37213 14139 37247
rect 16221 37213 16255 37247
rect 16313 37213 16347 37247
rect 16497 37213 16531 37247
rect 16584 37213 16618 37247
rect 17877 37213 17911 37247
rect 17969 37213 18003 37247
rect 18153 37213 18187 37247
rect 18245 37213 18279 37247
rect 20913 37213 20947 37247
rect 21281 37213 21315 37247
rect 25421 37213 25455 37247
rect 27261 37213 27295 37247
rect 9220 37145 9254 37179
rect 13001 37145 13035 37179
rect 14372 37145 14406 37179
rect 21097 37145 21131 37179
rect 21189 37145 21223 37179
rect 24777 37145 24811 37179
rect 25688 37145 25722 37179
rect 10333 37077 10367 37111
rect 12081 37077 12115 37111
rect 12265 37077 12299 37111
rect 13461 37077 13495 37111
rect 15485 37077 15519 37111
rect 21465 37077 21499 37111
rect 23673 37077 23707 37111
rect 23857 37077 23891 37111
rect 26801 37077 26835 37111
rect 11897 36873 11931 36907
rect 13461 36873 13495 36907
rect 14105 36873 14139 36907
rect 17049 36873 17083 36907
rect 18705 36873 18739 36907
rect 23121 36873 23155 36907
rect 23765 36873 23799 36907
rect 26433 36873 26467 36907
rect 27629 36873 27663 36907
rect 15761 36805 15795 36839
rect 19165 36805 19199 36839
rect 19365 36805 19399 36839
rect 28641 36805 28675 36839
rect 9597 36737 9631 36771
rect 9864 36737 9898 36771
rect 11713 36737 11747 36771
rect 11897 36737 11931 36771
rect 12357 36737 12391 36771
rect 12541 36737 12575 36771
rect 13369 36737 13403 36771
rect 13553 36737 13587 36771
rect 14013 36737 14047 36771
rect 14197 36737 14231 36771
rect 15577 36737 15611 36771
rect 15853 36737 15887 36771
rect 15945 36737 15979 36771
rect 16865 36737 16899 36771
rect 20361 36737 20395 36771
rect 20453 36737 20487 36771
rect 20637 36737 20671 36771
rect 20729 36737 20763 36771
rect 21833 36737 21867 36771
rect 22017 36737 22051 36771
rect 22109 36737 22143 36771
rect 22201 36737 22235 36771
rect 23029 36737 23063 36771
rect 23213 36737 23247 36771
rect 23673 36737 23707 36771
rect 23857 36737 23891 36771
rect 24501 36737 24535 36771
rect 25053 36737 25087 36771
rect 25320 36737 25354 36771
rect 27813 36737 27847 36771
rect 16681 36669 16715 36703
rect 18245 36669 18279 36703
rect 28273 36669 28307 36703
rect 12357 36601 12391 36635
rect 18613 36601 18647 36635
rect 28825 36601 28859 36635
rect 10977 36533 11011 36567
rect 16129 36533 16163 36567
rect 19349 36533 19383 36567
rect 19533 36533 19567 36567
rect 20177 36533 20211 36567
rect 22385 36533 22419 36567
rect 24317 36533 24351 36567
rect 28641 36533 28675 36567
rect 13185 36329 13219 36363
rect 16221 36329 16255 36363
rect 16957 36329 16991 36363
rect 18245 36329 18279 36363
rect 19625 36329 19659 36363
rect 22293 36329 22327 36363
rect 25697 36329 25731 36363
rect 19809 36261 19843 36295
rect 26341 36261 26375 36295
rect 17877 36193 17911 36227
rect 28549 36193 28583 36227
rect 11805 36125 11839 36159
rect 13185 36125 13219 36159
rect 13369 36125 13403 36159
rect 18061 36125 18095 36159
rect 19257 36125 19291 36159
rect 21005 36125 21039 36159
rect 21097 36125 21131 36159
rect 21281 36125 21315 36159
rect 21373 36125 21407 36159
rect 26525 36125 26559 36159
rect 28457 36125 28491 36159
rect 28641 36125 28675 36159
rect 16129 36057 16163 36091
rect 16865 36057 16899 36091
rect 19625 36057 19659 36091
rect 22109 36057 22143 36091
rect 25513 36057 25547 36091
rect 11621 35989 11655 36023
rect 20821 35989 20855 36023
rect 22309 35989 22343 36023
rect 22477 35989 22511 36023
rect 25713 35989 25747 36023
rect 25881 35989 25915 36023
rect 13553 35785 13587 35819
rect 26065 35785 26099 35819
rect 28115 35785 28149 35819
rect 28825 35785 28859 35819
rect 29745 35785 29779 35819
rect 10057 35717 10091 35751
rect 16948 35717 16982 35751
rect 22293 35717 22327 35751
rect 25881 35717 25915 35751
rect 27905 35717 27939 35751
rect 30389 35717 30423 35751
rect 30589 35717 30623 35751
rect 9873 35649 9907 35683
rect 11529 35649 11563 35683
rect 11785 35649 11819 35683
rect 13369 35649 13403 35683
rect 15485 35649 15519 35683
rect 15577 35649 15611 35683
rect 15761 35649 15795 35683
rect 15853 35649 15887 35683
rect 16681 35649 16715 35683
rect 19073 35649 19107 35683
rect 19901 35649 19935 35683
rect 20545 35649 20579 35683
rect 20729 35649 20763 35683
rect 23121 35649 23155 35683
rect 23388 35649 23422 35683
rect 28733 35649 28767 35683
rect 28917 35649 28951 35683
rect 29561 35649 29595 35683
rect 19717 35581 19751 35615
rect 20637 35581 20671 35615
rect 19257 35513 19291 35547
rect 21925 35513 21959 35547
rect 25513 35513 25547 35547
rect 10241 35445 10275 35479
rect 12909 35445 12943 35479
rect 15301 35445 15335 35479
rect 18061 35445 18095 35479
rect 20085 35445 20119 35479
rect 22293 35445 22327 35479
rect 22477 35445 22511 35479
rect 24501 35445 24535 35479
rect 25881 35445 25915 35479
rect 28089 35445 28123 35479
rect 28273 35445 28307 35479
rect 30573 35445 30607 35479
rect 30757 35445 30791 35479
rect 9873 35241 9907 35275
rect 11805 35241 11839 35275
rect 16773 35241 16807 35275
rect 17969 35241 18003 35275
rect 19257 35241 19291 35275
rect 21833 35241 21867 35275
rect 22293 35241 22327 35275
rect 23673 35241 23707 35275
rect 28181 35241 28215 35275
rect 30389 35241 30423 35275
rect 31033 35241 31067 35275
rect 12725 35173 12759 35207
rect 21649 35173 21683 35207
rect 25421 35173 25455 35207
rect 25973 35173 26007 35207
rect 30205 35173 30239 35207
rect 31217 35173 31251 35207
rect 11345 35105 11379 35139
rect 15301 35105 15335 35139
rect 15945 35105 15979 35139
rect 10149 35037 10183 35071
rect 10241 35037 10275 35071
rect 10333 35037 10367 35071
rect 10517 35037 10551 35071
rect 10977 35037 11011 35071
rect 11161 35037 11195 35071
rect 11805 35037 11839 35071
rect 11989 35037 12023 35071
rect 12541 35037 12575 35071
rect 14105 35037 14139 35071
rect 14198 35037 14232 35071
rect 14611 35037 14645 35071
rect 15485 35037 15519 35071
rect 15669 35037 15703 35071
rect 16405 35037 16439 35071
rect 16589 35037 16623 35071
rect 17969 35037 18003 35071
rect 18153 35037 18187 35071
rect 19257 35037 19291 35071
rect 19441 35037 19475 35071
rect 20729 35037 20763 35071
rect 20913 35037 20947 35071
rect 22477 35037 22511 35071
rect 25973 35037 26007 35071
rect 26157 35037 26191 35071
rect 27813 35037 27847 35071
rect 28825 35037 28859 35071
rect 29009 35037 29043 35071
rect 29929 35037 29963 35071
rect 14381 34969 14415 35003
rect 14473 34969 14507 35003
rect 15577 34969 15611 35003
rect 15807 34969 15841 35003
rect 20821 34969 20855 35003
rect 21373 34969 21407 35003
rect 23489 34969 23523 35003
rect 23705 34969 23739 35003
rect 25053 34969 25087 35003
rect 28181 34969 28215 35003
rect 28917 34969 28951 35003
rect 30849 34969 30883 35003
rect 14749 34901 14783 34935
rect 23857 34901 23891 34935
rect 25513 34901 25547 34935
rect 28365 34901 28399 34935
rect 31059 34901 31093 34935
rect 8677 34697 8711 34731
rect 12725 34697 12759 34731
rect 14289 34697 14323 34731
rect 21189 34697 21223 34731
rect 22201 34697 22235 34731
rect 22753 34697 22787 34731
rect 23857 34697 23891 34731
rect 25789 34697 25823 34731
rect 27997 34697 28031 34731
rect 29745 34697 29779 34731
rect 31585 34697 31619 34731
rect 12449 34629 12483 34663
rect 17049 34629 17083 34663
rect 18981 34629 19015 34663
rect 19073 34629 19107 34663
rect 19191 34629 19225 34663
rect 20177 34629 20211 34663
rect 20407 34629 20441 34663
rect 8953 34561 8987 34595
rect 9045 34561 9079 34595
rect 9137 34561 9171 34595
rect 9321 34561 9355 34595
rect 12081 34561 12115 34595
rect 12229 34561 12263 34595
rect 12357 34561 12391 34595
rect 12587 34561 12621 34595
rect 13645 34561 13679 34595
rect 13793 34561 13827 34595
rect 13921 34561 13955 34595
rect 14013 34561 14047 34595
rect 14151 34561 14185 34595
rect 15485 34561 15519 34595
rect 16865 34561 16899 34595
rect 16957 34561 16991 34595
rect 17167 34561 17201 34595
rect 17325 34561 17359 34595
rect 18889 34561 18923 34595
rect 20085 34561 20119 34595
rect 20269 34561 20303 34595
rect 21097 34561 21131 34595
rect 21281 34561 21315 34595
rect 22017 34561 22051 34595
rect 22661 34561 22695 34595
rect 22820 34561 22854 34595
rect 25697 34561 25731 34595
rect 25881 34561 25915 34595
rect 28457 34561 28491 34595
rect 28641 34561 28675 34595
rect 30205 34561 30239 34595
rect 30472 34561 30506 34595
rect 9781 34493 9815 34527
rect 10057 34493 10091 34527
rect 15209 34493 15243 34527
rect 19349 34493 19383 34527
rect 20545 34493 20579 34527
rect 21833 34493 21867 34527
rect 23397 34493 23431 34527
rect 27537 34493 27571 34527
rect 29285 34493 29319 34527
rect 23673 34425 23707 34459
rect 27813 34425 27847 34459
rect 28457 34425 28491 34459
rect 29653 34425 29687 34459
rect 16681 34357 16715 34391
rect 18705 34357 18739 34391
rect 19901 34357 19935 34391
rect 9413 34153 9447 34187
rect 16865 34153 16899 34187
rect 23673 34153 23707 34187
rect 30573 34153 30607 34187
rect 31217 34153 31251 34187
rect 13369 34085 13403 34119
rect 29561 34085 29595 34119
rect 30205 34085 30239 34119
rect 10793 34017 10827 34051
rect 9689 33949 9723 33983
rect 9781 33949 9815 33983
rect 9873 33949 9907 33983
rect 10057 33949 10091 33983
rect 10517 33949 10551 33983
rect 12173 33949 12207 33983
rect 12321 33949 12355 33983
rect 12449 33949 12483 33983
rect 12679 33949 12713 33983
rect 13553 33949 13587 33983
rect 14933 33949 14967 33983
rect 15209 33949 15243 33983
rect 16221 33949 16255 33983
rect 16314 33949 16348 33983
rect 16497 33949 16531 33983
rect 16589 33949 16623 33983
rect 16686 33949 16720 33983
rect 17417 33949 17451 33983
rect 17693 33949 17727 33983
rect 19257 33949 19291 33983
rect 19405 33949 19439 33983
rect 19761 33949 19795 33983
rect 20453 33949 20487 33983
rect 20546 33949 20580 33983
rect 20821 33949 20855 33983
rect 20959 33949 20993 33983
rect 21649 33949 21683 33983
rect 21797 33949 21831 33983
rect 22017 33949 22051 33983
rect 22114 33949 22148 33983
rect 23305 33949 23339 33983
rect 24593 33949 24627 33983
rect 28089 33949 28123 33983
rect 29561 33949 29595 33983
rect 29745 33949 29779 33983
rect 31401 33949 31435 33983
rect 12541 33881 12575 33915
rect 19533 33881 19567 33915
rect 19645 33881 19679 33915
rect 20729 33881 20763 33915
rect 21925 33881 21959 33915
rect 25697 33881 25731 33915
rect 12817 33813 12851 33847
rect 19901 33813 19935 33847
rect 21097 33813 21131 33847
rect 22293 33813 22327 33847
rect 23673 33813 23707 33847
rect 23857 33813 23891 33847
rect 24409 33813 24443 33847
rect 26985 33813 27019 33847
rect 27905 33813 27939 33847
rect 30573 33813 30607 33847
rect 30757 33813 30791 33847
rect 10425 33609 10459 33643
rect 11989 33609 12023 33643
rect 13645 33609 13679 33643
rect 15945 33609 15979 33643
rect 20545 33609 20579 33643
rect 24225 33609 24259 33643
rect 26433 33609 26467 33643
rect 29561 33609 29595 33643
rect 10057 33541 10091 33575
rect 12357 33541 12391 33575
rect 12475 33541 12509 33575
rect 14151 33541 14185 33575
rect 20821 33541 20855 33575
rect 20913 33541 20947 33575
rect 25320 33541 25354 33575
rect 30297 33541 30331 33575
rect 10241 33473 10275 33507
rect 12173 33473 12207 33507
rect 12265 33473 12299 33507
rect 13829 33473 13863 33507
rect 13921 33473 13955 33507
rect 14013 33473 14047 33507
rect 14933 33473 14967 33507
rect 15025 33473 15059 33507
rect 15117 33473 15151 33507
rect 15255 33473 15289 33507
rect 15853 33473 15887 33507
rect 16037 33473 16071 33507
rect 18245 33473 18279 33507
rect 20729 33473 20763 33507
rect 21031 33473 21065 33507
rect 22457 33473 22491 33507
rect 24133 33473 24167 33507
rect 24317 33473 24351 33507
rect 25053 33473 25087 33507
rect 27537 33473 27571 33507
rect 27804 33473 27838 33507
rect 29469 33473 29503 33507
rect 30205 33473 30239 33507
rect 30389 33473 30423 33507
rect 12633 33405 12667 33439
rect 14289 33405 14323 33439
rect 15393 33405 15427 33439
rect 16681 33405 16715 33439
rect 16957 33405 16991 33439
rect 17969 33405 18003 33439
rect 19257 33405 19291 33439
rect 21189 33405 21223 33439
rect 22201 33405 22235 33439
rect 19487 33337 19521 33371
rect 14749 33269 14783 33303
rect 23581 33269 23615 33303
rect 28917 33269 28951 33303
rect 21925 33065 21959 33099
rect 29009 33065 29043 33099
rect 12081 32997 12115 33031
rect 20453 32997 20487 33031
rect 11161 32929 11195 32963
rect 14105 32929 14139 32963
rect 16221 32929 16255 32963
rect 17877 32929 17911 32963
rect 9045 32861 9079 32895
rect 9965 32861 9999 32895
rect 10054 32861 10088 32895
rect 10149 32861 10183 32895
rect 10333 32861 10367 32895
rect 10793 32861 10827 32895
rect 10977 32861 11011 32895
rect 12265 32861 12299 32895
rect 12357 32861 12391 32895
rect 12725 32861 12759 32895
rect 16497 32861 16531 32895
rect 17601 32861 17635 32895
rect 19257 32861 19291 32895
rect 19441 32861 19475 32895
rect 19625 32861 19659 32895
rect 19717 32861 19751 32895
rect 22109 32861 22143 32895
rect 22385 32861 22419 32895
rect 24961 32861 24995 32895
rect 27629 32861 27663 32895
rect 30757 32861 30791 32895
rect 9229 32793 9263 32827
rect 12449 32793 12483 32827
rect 12587 32793 12621 32827
rect 14372 32793 14406 32827
rect 20269 32793 20303 32827
rect 23397 32793 23431 32827
rect 23581 32793 23615 32827
rect 25228 32793 25262 32827
rect 27896 32793 27930 32827
rect 9689 32725 9723 32759
rect 15485 32725 15519 32759
rect 22293 32725 22327 32759
rect 26341 32725 26375 32759
rect 30573 32725 30607 32759
rect 10977 32521 11011 32555
rect 16037 32521 16071 32555
rect 20453 32521 20487 32555
rect 22477 32521 22511 32555
rect 24501 32521 24535 32555
rect 25329 32521 25363 32555
rect 28181 32521 28215 32555
rect 28549 32521 28583 32555
rect 31585 32521 31619 32555
rect 9842 32453 9876 32487
rect 11529 32453 11563 32487
rect 14933 32453 14967 32487
rect 15025 32453 15059 32487
rect 17049 32453 17083 32487
rect 18696 32453 18730 32487
rect 30472 32453 30506 32487
rect 5825 32385 5859 32419
rect 6561 32385 6595 32419
rect 7941 32385 7975 32419
rect 11713 32385 11747 32419
rect 13461 32385 13495 32419
rect 14657 32385 14691 32419
rect 14805 32385 14839 32419
rect 15122 32385 15156 32419
rect 15945 32385 15979 32419
rect 16773 32385 16807 32419
rect 16921 32385 16955 32419
rect 17141 32385 17175 32419
rect 17279 32385 17313 32419
rect 20361 32385 20395 32419
rect 24409 32385 24443 32419
rect 24593 32385 24627 32419
rect 25513 32385 25547 32419
rect 25697 32385 25731 32419
rect 25789 32385 25823 32419
rect 27445 32385 27479 32419
rect 27629 32385 27663 32419
rect 27721 32385 27755 32419
rect 28365 32385 28399 32419
rect 28641 32385 28675 32419
rect 9597 32317 9631 32351
rect 13001 32317 13035 32351
rect 13369 32317 13403 32351
rect 18429 32317 18463 32351
rect 21833 32317 21867 32351
rect 22201 32317 22235 32351
rect 22293 32317 22327 32351
rect 30205 32317 30239 32351
rect 19809 32249 19843 32283
rect 5641 32181 5675 32215
rect 6377 32181 6411 32215
rect 7757 32181 7791 32215
rect 11897 32181 11931 32215
rect 13645 32181 13679 32215
rect 15301 32181 15335 32215
rect 17417 32181 17451 32215
rect 27261 32181 27295 32215
rect 10609 31977 10643 32011
rect 13553 31977 13587 32011
rect 16957 31977 16991 32011
rect 19901 31977 19935 32011
rect 26065 31977 26099 32011
rect 28089 31977 28123 32011
rect 30481 31977 30515 32011
rect 30665 31977 30699 32011
rect 17877 31909 17911 31943
rect 22017 31909 22051 31943
rect 30113 31909 30147 31943
rect 31125 31909 31159 31943
rect 19257 31841 19291 31875
rect 22477 31841 22511 31875
rect 25881 31841 25915 31875
rect 27813 31841 27847 31875
rect 4997 31773 5031 31807
rect 7021 31773 7055 31807
rect 7288 31773 7322 31807
rect 9229 31773 9263 31807
rect 12173 31773 12207 31807
rect 12440 31773 12474 31807
rect 14105 31773 14139 31807
rect 14289 31773 14323 31807
rect 14473 31773 14507 31807
rect 14565 31773 14599 31807
rect 15669 31773 15703 31807
rect 18061 31773 18095 31807
rect 18153 31773 18187 31807
rect 18245 31773 18279 31807
rect 18363 31773 18397 31807
rect 18521 31773 18555 31807
rect 19625 31773 19659 31807
rect 19717 31773 19751 31807
rect 20637 31773 20671 31807
rect 25789 31773 25823 31807
rect 27905 31773 27939 31807
rect 31125 31773 31159 31807
rect 31309 31773 31343 31807
rect 5264 31705 5298 31739
rect 9496 31705 9530 31739
rect 20904 31705 20938 31739
rect 22744 31705 22778 31739
rect 6377 31637 6411 31671
rect 8401 31637 8435 31671
rect 23857 31637 23891 31671
rect 25421 31637 25455 31671
rect 27445 31637 27479 31671
rect 30481 31637 30515 31671
rect 5825 31433 5859 31467
rect 6577 31433 6611 31467
rect 6745 31433 6779 31467
rect 9597 31433 9631 31467
rect 12909 31433 12943 31467
rect 13737 31433 13771 31467
rect 20821 31433 20855 31467
rect 21189 31433 21223 31467
rect 21833 31433 21867 31467
rect 27537 31433 27571 31467
rect 28181 31433 28215 31467
rect 30849 31433 30883 31467
rect 5457 31365 5491 31399
rect 5673 31365 5707 31399
rect 6377 31365 6411 31399
rect 16681 31365 16715 31399
rect 19073 31365 19107 31399
rect 19257 31365 19291 31399
rect 22477 31365 22511 31399
rect 23213 31365 23247 31399
rect 7205 31297 7239 31331
rect 7461 31297 7495 31331
rect 9873 31297 9907 31331
rect 9965 31297 9999 31331
rect 10057 31297 10091 31331
rect 10241 31297 10275 31331
rect 11529 31297 11563 31331
rect 11796 31297 11830 31331
rect 13369 31297 13403 31331
rect 13553 31297 13587 31331
rect 13829 31297 13863 31331
rect 14289 31297 14323 31331
rect 14545 31297 14579 31331
rect 16865 31297 16899 31331
rect 18153 31297 18187 31331
rect 20177 31297 20211 31331
rect 21005 31297 21039 31331
rect 21281 31297 21315 31331
rect 22293 31297 22327 31331
rect 23673 31297 23707 31331
rect 24961 31297 24995 31331
rect 25228 31297 25262 31331
rect 27997 31297 28031 31331
rect 28917 31297 28951 31331
rect 29184 31297 29218 31331
rect 30757 31297 30791 31331
rect 30941 31297 30975 31331
rect 22201 31229 22235 31263
rect 23581 31229 23615 31263
rect 27905 31229 27939 31263
rect 18337 31161 18371 31195
rect 5641 31093 5675 31127
rect 6561 31093 6595 31127
rect 8585 31093 8619 31127
rect 15669 31093 15703 31127
rect 17049 31093 17083 31127
rect 20269 31093 20303 31127
rect 23857 31093 23891 31127
rect 26341 31093 26375 31127
rect 30297 31093 30331 31127
rect 6377 30889 6411 30923
rect 7113 30889 7147 30923
rect 7941 30889 7975 30923
rect 8125 30889 8159 30923
rect 12725 30889 12759 30923
rect 14105 30889 14139 30923
rect 23121 30889 23155 30923
rect 24501 30889 24535 30923
rect 18705 30821 18739 30855
rect 4997 30753 5031 30787
rect 12081 30753 12115 30787
rect 12449 30753 12483 30787
rect 15485 30753 15519 30787
rect 17325 30753 17359 30787
rect 19625 30753 19659 30787
rect 25789 30753 25823 30787
rect 28273 30753 28307 30787
rect 5264 30685 5298 30719
rect 7297 30685 7331 30719
rect 12541 30685 12575 30719
rect 14381 30685 14415 30719
rect 14473 30685 14507 30719
rect 14565 30685 14599 30719
rect 14749 30685 14783 30719
rect 19717 30685 19751 30719
rect 23305 30685 23339 30719
rect 23581 30685 23615 30719
rect 24685 30685 24719 30719
rect 24869 30685 24903 30719
rect 24961 30685 24995 30719
rect 25881 30685 25915 30719
rect 28181 30685 28215 30719
rect 7757 30617 7791 30651
rect 15752 30617 15786 30651
rect 17592 30617 17626 30651
rect 19257 30617 19291 30651
rect 26065 30617 26099 30651
rect 7957 30549 7991 30583
rect 16865 30549 16899 30583
rect 19901 30549 19935 30583
rect 23489 30549 23523 30583
rect 25421 30549 25455 30583
rect 27813 30549 27847 30583
rect 28457 30549 28491 30583
rect 8125 30345 8159 30379
rect 17785 30345 17819 30379
rect 18797 30345 18831 30379
rect 22661 30345 22695 30379
rect 24593 30345 24627 30379
rect 28273 30345 28307 30379
rect 7757 30277 7791 30311
rect 7973 30277 8007 30311
rect 13645 30277 13679 30311
rect 15209 30277 15243 30311
rect 16681 30277 16715 30311
rect 20637 30277 20671 30311
rect 25973 30277 26007 30311
rect 27905 30277 27939 30311
rect 13461 30209 13495 30243
rect 14841 30209 14875 30243
rect 15025 30209 15059 30243
rect 16957 30209 16991 30243
rect 17049 30209 17083 30243
rect 17141 30209 17175 30243
rect 17325 30209 17359 30243
rect 17969 30209 18003 30243
rect 18153 30209 18187 30243
rect 18245 30209 18279 30243
rect 18705 30209 18739 30243
rect 18889 30209 18923 30243
rect 20453 30209 20487 30243
rect 22569 30209 22603 30243
rect 23469 30209 23503 30243
rect 28089 30209 28123 30243
rect 28349 30199 28383 30233
rect 23213 30141 23247 30175
rect 7941 30005 7975 30039
rect 26065 30005 26099 30039
rect 5641 29801 5675 29835
rect 9505 29801 9539 29835
rect 11529 29801 11563 29835
rect 18613 29801 18647 29835
rect 22109 29801 22143 29835
rect 23121 29801 23155 29835
rect 26801 29801 26835 29835
rect 28917 29801 28951 29835
rect 33333 29801 33367 29835
rect 31493 29733 31527 29767
rect 27537 29665 27571 29699
rect 4997 29597 5031 29631
rect 6469 29597 6503 29631
rect 7941 29597 7975 29631
rect 10149 29597 10183 29631
rect 11989 29597 12023 29631
rect 12817 29597 12851 29631
rect 14289 29597 14323 29631
rect 23351 29597 23385 29631
rect 23470 29597 23504 29631
rect 23581 29597 23615 29631
rect 23765 29597 23799 29631
rect 24409 29597 24443 29631
rect 25421 29597 25455 29631
rect 30113 29597 30147 29631
rect 31953 29597 31987 29631
rect 5457 29529 5491 29563
rect 5673 29529 5707 29563
rect 9321 29529 9355 29563
rect 10416 29529 10450 29563
rect 12173 29529 12207 29563
rect 13001 29529 13035 29563
rect 14105 29529 14139 29563
rect 18521 29529 18555 29563
rect 19257 29529 19291 29563
rect 19441 29529 19475 29563
rect 20637 29529 20671 29563
rect 25688 29529 25722 29563
rect 27804 29529 27838 29563
rect 30358 29529 30392 29563
rect 32198 29529 32232 29563
rect 4813 29461 4847 29495
rect 5825 29461 5859 29495
rect 6285 29461 6319 29495
rect 7757 29461 7791 29495
rect 9521 29461 9555 29495
rect 9689 29461 9723 29495
rect 12357 29461 12391 29495
rect 13185 29461 13219 29495
rect 14473 29461 14507 29495
rect 19625 29461 19659 29495
rect 24593 29461 24627 29495
rect 10425 29257 10459 29291
rect 11621 29257 11655 29291
rect 14105 29257 14139 29291
rect 15945 29257 15979 29291
rect 23213 29257 23247 29291
rect 24041 29257 24075 29291
rect 25421 29257 25455 29291
rect 27721 29257 27755 29291
rect 29653 29257 29687 29291
rect 4712 29189 4746 29223
rect 6377 29189 6411 29223
rect 6577 29189 6611 29223
rect 24777 29189 24811 29223
rect 4445 29121 4479 29155
rect 8033 29121 8067 29155
rect 9045 29121 9079 29155
rect 9312 29121 9346 29155
rect 11897 29121 11931 29155
rect 11989 29121 12023 29155
rect 12081 29121 12115 29155
rect 12265 29121 12299 29155
rect 12725 29121 12759 29155
rect 12981 29121 13015 29155
rect 14565 29121 14599 29155
rect 14821 29121 14855 29155
rect 17877 29121 17911 29155
rect 19257 29121 19291 29155
rect 19524 29121 19558 29155
rect 21833 29121 21867 29155
rect 22100 29121 22134 29155
rect 23673 29121 23707 29155
rect 23857 29121 23891 29155
rect 24593 29121 24627 29155
rect 25651 29121 25685 29155
rect 25789 29121 25823 29155
rect 25881 29121 25915 29155
rect 26065 29121 26099 29155
rect 28825 29121 28859 29155
rect 29009 29121 29043 29155
rect 29929 29121 29963 29155
rect 30021 29121 30055 29155
rect 30113 29121 30147 29155
rect 30297 29121 30331 29155
rect 7757 29053 7791 29087
rect 17693 29053 17727 29087
rect 28089 29053 28123 29087
rect 28181 29053 28215 29087
rect 5825 28985 5859 29019
rect 6745 28985 6779 29019
rect 18061 28985 18095 29019
rect 20637 28985 20671 29019
rect 29193 28985 29227 29019
rect 6561 28917 6595 28951
rect 28365 28917 28399 28951
rect 6837 28713 6871 28747
rect 7941 28713 7975 28747
rect 12725 28713 12759 28747
rect 14565 28713 14599 28747
rect 20729 28713 20763 28747
rect 21833 28713 21867 28747
rect 24593 28713 24627 28747
rect 25697 28713 25731 28747
rect 27629 28713 27663 28747
rect 29745 28713 29779 28747
rect 32413 28713 32447 28747
rect 8125 28645 8159 28679
rect 18613 28645 18647 28679
rect 28825 28645 28859 28679
rect 15761 28577 15795 28611
rect 23305 28577 23339 28611
rect 5549 28509 5583 28543
rect 10517 28509 10551 28543
rect 13001 28509 13035 28543
rect 13093 28509 13127 28543
rect 13185 28509 13219 28543
rect 13369 28509 13403 28543
rect 14841 28509 14875 28543
rect 14930 28509 14964 28543
rect 15030 28509 15064 28543
rect 15209 28509 15243 28543
rect 18061 28509 18095 28543
rect 18429 28509 18463 28543
rect 19717 28509 19751 28543
rect 19901 28509 19935 28543
rect 19993 28509 20027 28543
rect 20177 28509 20211 28543
rect 20269 28509 20303 28543
rect 21005 28509 21039 28543
rect 21097 28509 21131 28543
rect 21189 28509 21223 28543
rect 21373 28509 21407 28543
rect 22063 28509 22097 28543
rect 22201 28509 22235 28543
rect 22293 28509 22327 28543
rect 22477 28509 22511 28543
rect 25329 28509 25363 28543
rect 27813 28509 27847 28543
rect 28089 28509 28123 28543
rect 30021 28509 30055 28543
rect 30113 28509 30147 28543
rect 30205 28509 30239 28543
rect 30389 28509 30423 28543
rect 7757 28441 7791 28475
rect 7957 28441 7991 28475
rect 16006 28441 16040 28475
rect 18245 28441 18279 28475
rect 18337 28441 18371 28475
rect 22937 28441 22971 28475
rect 23121 28441 23155 28475
rect 24409 28441 24443 28475
rect 25513 28441 25547 28475
rect 26985 28441 27019 28475
rect 28641 28441 28675 28475
rect 31125 28441 31159 28475
rect 11805 28373 11839 28407
rect 17141 28373 17175 28407
rect 24609 28373 24643 28407
rect 24777 28373 24811 28407
rect 27077 28373 27111 28407
rect 27997 28373 28031 28407
rect 6653 28169 6687 28203
rect 8677 28169 8711 28203
rect 13645 28169 13679 28203
rect 15485 28169 15519 28203
rect 18245 28169 18279 28203
rect 19073 28169 19107 28203
rect 21189 28169 21223 28203
rect 26433 28169 26467 28203
rect 31033 28169 31067 28203
rect 19901 28101 19935 28135
rect 24225 28101 24259 28135
rect 27353 28101 27387 28135
rect 6837 28033 6871 28067
rect 7297 28033 7331 28067
rect 7564 28033 7598 28067
rect 9137 28033 9171 28067
rect 9393 28033 9427 28067
rect 11529 28033 11563 28067
rect 11785 28033 11819 28067
rect 13553 28033 13587 28067
rect 14841 28033 14875 28067
rect 15761 28033 15795 28067
rect 15853 28033 15887 28067
rect 15966 28033 16000 28067
rect 16129 28033 16163 28067
rect 16865 28033 16899 28067
rect 17132 28033 17166 28067
rect 18889 28033 18923 28067
rect 19717 28033 19751 28067
rect 21005 28033 21039 28067
rect 21925 28033 21959 28067
rect 22192 28033 22226 28067
rect 25053 28033 25087 28067
rect 25320 28033 25354 28067
rect 29791 28033 29825 28067
rect 29929 28033 29963 28067
rect 30021 28036 30055 28070
rect 30205 28033 30239 28067
rect 30665 28033 30699 28067
rect 30849 28033 30883 28067
rect 20821 27965 20855 27999
rect 12909 27897 12943 27931
rect 23305 27897 23339 27931
rect 23857 27897 23891 27931
rect 10517 27829 10551 27863
rect 14933 27829 14967 27863
rect 24225 27829 24259 27863
rect 24409 27829 24443 27863
rect 28641 27829 28675 27863
rect 29561 27829 29595 27863
rect 6745 27625 6779 27659
rect 7941 27625 7975 27659
rect 11253 27625 11287 27659
rect 17509 27625 17543 27659
rect 10701 27557 10735 27591
rect 16773 27557 16807 27591
rect 21557 27557 21591 27591
rect 24685 27557 24719 27591
rect 26433 27557 26467 27591
rect 12817 27489 12851 27523
rect 21097 27489 21131 27523
rect 5365 27421 5399 27455
rect 5632 27421 5666 27455
rect 10517 27421 10551 27455
rect 11529 27421 11563 27455
rect 11621 27421 11655 27455
rect 11713 27421 11747 27455
rect 11897 27421 11931 27455
rect 12633 27421 12667 27455
rect 13277 27421 13311 27455
rect 15393 27421 15427 27455
rect 17693 27421 17727 27455
rect 19533 27421 19567 27455
rect 19625 27421 19659 27455
rect 19717 27421 19751 27455
rect 19901 27421 19935 27455
rect 20913 27421 20947 27455
rect 21833 27421 21867 27455
rect 21925 27421 21959 27455
rect 22017 27421 22051 27455
rect 22201 27421 22235 27455
rect 22845 27421 22879 27455
rect 25789 27421 25823 27455
rect 25882 27421 25916 27455
rect 26157 27421 26191 27455
rect 26254 27421 26288 27455
rect 27077 27421 27111 27455
rect 27813 27421 27847 27455
rect 27961 27421 27995 27455
rect 28278 27421 28312 27455
rect 29837 27421 29871 27455
rect 29929 27421 29963 27455
rect 30021 27421 30055 27455
rect 30205 27421 30239 27455
rect 7757 27353 7791 27387
rect 7957 27353 7991 27387
rect 12449 27353 12483 27387
rect 14565 27353 14599 27387
rect 14749 27353 14783 27387
rect 15638 27353 15672 27387
rect 20729 27353 20763 27387
rect 23673 27353 23707 27387
rect 24409 27353 24443 27387
rect 26065 27353 26099 27387
rect 26893 27353 26927 27387
rect 28089 27353 28123 27387
rect 28181 27353 28215 27387
rect 8125 27285 8159 27319
rect 13461 27285 13495 27319
rect 14933 27285 14967 27319
rect 19257 27285 19291 27319
rect 23029 27285 23063 27319
rect 23765 27285 23799 27319
rect 24869 27285 24903 27319
rect 27261 27285 27295 27319
rect 28457 27285 28491 27319
rect 29561 27285 29595 27319
rect 7205 27081 7239 27115
rect 7849 27081 7883 27115
rect 10425 27081 10459 27115
rect 15393 27081 15427 27115
rect 17233 27081 17267 27115
rect 24133 27081 24167 27115
rect 24777 27081 24811 27115
rect 25421 27081 25455 27115
rect 28089 27081 28123 27115
rect 31217 27081 31251 27115
rect 6377 27013 6411 27047
rect 6577 27013 6611 27047
rect 22477 27013 22511 27047
rect 23213 27013 23247 27047
rect 27721 27013 27755 27047
rect 28917 27013 28951 27047
rect 30082 27013 30116 27047
rect 4445 26945 4479 26979
rect 4712 26945 4746 26979
rect 7389 26945 7423 26979
rect 8033 26945 8067 26979
rect 8677 26945 8711 26979
rect 9965 26945 9999 26979
rect 10609 26945 10643 26979
rect 13921 26945 13955 26979
rect 15669 26945 15703 26979
rect 15761 26945 15795 26979
rect 15853 26945 15887 26979
rect 16037 26945 16071 26979
rect 17141 26945 17175 26979
rect 17969 26945 18003 26979
rect 18613 26945 18647 26979
rect 18880 26945 18914 26979
rect 21005 26945 21039 26979
rect 21189 26945 21223 26979
rect 21281 26945 21315 26979
rect 22293 26945 22327 26979
rect 23397 26945 23431 26979
rect 24041 26945 24075 26979
rect 24225 26945 24259 26979
rect 24685 26945 24719 26979
rect 24869 26945 24903 26979
rect 25697 26945 25731 26979
rect 25789 26945 25823 26979
rect 25881 26945 25915 26979
rect 26065 26945 26099 26979
rect 27077 26945 27111 26979
rect 27905 26945 27939 26979
rect 28549 26945 28583 26979
rect 28697 26945 28731 26979
rect 28825 26945 28859 26979
rect 29014 26945 29048 26979
rect 13553 26877 13587 26911
rect 14013 26877 14047 26911
rect 18153 26877 18187 26911
rect 21833 26877 21867 26911
rect 22201 26877 22235 26911
rect 29837 26877 29871 26911
rect 19993 26809 20027 26843
rect 27261 26809 27295 26843
rect 5825 26741 5859 26775
rect 6561 26741 6595 26775
rect 6745 26741 6779 26775
rect 8493 26741 8527 26775
rect 9781 26741 9815 26775
rect 14197 26741 14231 26775
rect 20821 26741 20855 26775
rect 23581 26741 23615 26775
rect 29193 26741 29227 26775
rect 12633 26537 12667 26571
rect 15485 26537 15519 26571
rect 28825 26537 28859 26571
rect 31401 26537 31435 26571
rect 22017 26469 22051 26503
rect 11253 26401 11287 26435
rect 19533 26401 19567 26435
rect 20637 26401 20671 26435
rect 4905 26333 4939 26367
rect 7021 26333 7055 26367
rect 8953 26333 8987 26367
rect 13277 26333 13311 26367
rect 13461 26333 13495 26367
rect 13553 26333 13587 26367
rect 14105 26333 14139 26367
rect 19257 26333 19291 26367
rect 20904 26333 20938 26367
rect 22937 26333 22971 26367
rect 23029 26333 23063 26367
rect 23121 26333 23155 26367
rect 23305 26333 23339 26367
rect 28457 26333 28491 26367
rect 28641 26333 28675 26367
rect 30021 26333 30055 26367
rect 30288 26333 30322 26367
rect 5172 26265 5206 26299
rect 7288 26265 7322 26299
rect 9220 26265 9254 26299
rect 11520 26265 11554 26299
rect 13093 26265 13127 26299
rect 14350 26265 14384 26299
rect 6285 26197 6319 26231
rect 8401 26197 8435 26231
rect 10333 26197 10367 26231
rect 22661 26197 22695 26231
rect 5549 25993 5583 26027
rect 8125 25993 8159 26027
rect 10793 25993 10827 26027
rect 13645 25993 13679 26027
rect 14105 25993 14139 26027
rect 14473 25993 14507 26027
rect 15945 25993 15979 26027
rect 18245 25993 18279 26027
rect 19349 25993 19383 26027
rect 21097 25993 21131 26027
rect 25237 25993 25271 26027
rect 6377 25925 6411 25959
rect 6577 25925 6611 25959
rect 7757 25925 7791 25959
rect 7957 25925 7991 25959
rect 15577 25925 15611 25959
rect 18981 25925 19015 25959
rect 19165 25925 19199 25959
rect 20269 25925 20303 25959
rect 30481 25925 30515 25959
rect 5733 25857 5767 25891
rect 8953 25857 8987 25891
rect 9220 25857 9254 25891
rect 10977 25857 11011 25891
rect 13461 25857 13495 25891
rect 14289 25857 14323 25891
rect 14565 25857 14599 25891
rect 15761 25857 15795 25891
rect 16865 25857 16899 25891
rect 17132 25857 17166 25891
rect 21005 25857 21039 25891
rect 22661 25857 22695 25891
rect 25145 25857 25179 25891
rect 25329 25857 25363 25891
rect 25789 25857 25823 25891
rect 25882 25857 25916 25891
rect 26065 25857 26099 25891
rect 26157 25857 26191 25891
rect 26295 25857 26329 25891
rect 27241 25857 27275 25891
rect 30113 25857 30147 25891
rect 30206 25857 30240 25891
rect 30389 25857 30423 25891
rect 30619 25857 30653 25891
rect 13001 25789 13035 25823
rect 13369 25789 13403 25823
rect 26985 25789 27019 25823
rect 6745 25721 6779 25755
rect 6561 25653 6595 25687
rect 7941 25653 7975 25687
rect 10333 25653 10367 25687
rect 20361 25653 20395 25687
rect 22753 25653 22787 25687
rect 26433 25653 26467 25687
rect 28365 25653 28399 25687
rect 30757 25653 30791 25687
rect 5457 25449 5491 25483
rect 9137 25449 9171 25483
rect 10057 25449 10091 25483
rect 10241 25449 10275 25483
rect 10885 25449 10919 25483
rect 11989 25449 12023 25483
rect 17417 25449 17451 25483
rect 21373 25449 21407 25483
rect 26249 25449 26283 25483
rect 15209 25313 15243 25347
rect 5641 25245 5675 25279
rect 6929 25245 6963 25279
rect 8953 25245 8987 25279
rect 12817 25245 12851 25279
rect 15485 25245 15519 25279
rect 16773 25245 16807 25279
rect 17693 25245 17727 25279
rect 17785 25245 17819 25279
rect 17882 25242 17916 25276
rect 18061 25245 18095 25279
rect 19881 25245 19915 25279
rect 19993 25245 20027 25279
rect 20106 25245 20140 25279
rect 20269 25245 20303 25279
rect 21189 25245 21223 25279
rect 22477 25245 22511 25279
rect 22744 25245 22778 25279
rect 24409 25245 24443 25279
rect 26525 25245 26559 25279
rect 26614 25239 26648 25273
rect 26709 25245 26743 25279
rect 26893 25245 26927 25279
rect 27813 25245 27847 25279
rect 27906 25245 27940 25279
rect 28181 25245 28215 25279
rect 28319 25245 28353 25279
rect 30389 25245 30423 25279
rect 30537 25245 30571 25279
rect 30757 25245 30791 25279
rect 30854 25245 30888 25279
rect 9873 25177 9907 25211
rect 10701 25177 10735 25211
rect 11805 25177 11839 25211
rect 16589 25177 16623 25211
rect 19625 25177 19659 25211
rect 24654 25177 24688 25211
rect 28089 25177 28123 25211
rect 30665 25177 30699 25211
rect 6745 25109 6779 25143
rect 10073 25109 10107 25143
rect 10901 25109 10935 25143
rect 11069 25109 11103 25143
rect 12005 25109 12039 25143
rect 12173 25109 12207 25143
rect 12909 25109 12943 25143
rect 16957 25109 16991 25143
rect 23857 25109 23891 25143
rect 25789 25109 25823 25143
rect 28457 25109 28491 25143
rect 31033 25109 31067 25143
rect 9597 24905 9631 24939
rect 12909 24905 12943 24939
rect 21097 24905 21131 24939
rect 24041 24905 24075 24939
rect 26341 24905 26375 24939
rect 28365 24905 28399 24939
rect 29009 24905 29043 24939
rect 6929 24837 6963 24871
rect 7129 24837 7163 24871
rect 17877 24837 17911 24871
rect 19984 24837 20018 24871
rect 22753 24837 22787 24871
rect 4721 24769 4755 24803
rect 9781 24769 9815 24803
rect 10977 24769 11011 24803
rect 11785 24769 11819 24803
rect 13645 24769 13679 24803
rect 13737 24769 13771 24803
rect 13829 24769 13863 24803
rect 14013 24769 14047 24803
rect 14924 24769 14958 24803
rect 16957 24769 16991 24803
rect 17049 24769 17083 24803
rect 17141 24769 17175 24803
rect 17325 24769 17359 24803
rect 18061 24769 18095 24803
rect 18705 24769 18739 24803
rect 18889 24769 18923 24803
rect 19717 24769 19751 24803
rect 21925 24769 21959 24803
rect 24317 24769 24351 24803
rect 24409 24769 24443 24803
rect 24501 24769 24535 24803
rect 24685 24769 24719 24803
rect 25237 24769 25271 24803
rect 25973 24769 26007 24803
rect 26157 24769 26191 24803
rect 27241 24769 27275 24803
rect 28825 24769 28859 24803
rect 30389 24769 30423 24803
rect 30481 24769 30515 24803
rect 30573 24769 30607 24803
rect 30757 24769 30791 24803
rect 31217 24769 31251 24803
rect 31401 24769 31435 24803
rect 11529 24701 11563 24735
rect 14657 24701 14691 24735
rect 16681 24701 16715 24735
rect 18245 24701 18279 24735
rect 26985 24701 27019 24735
rect 10793 24633 10827 24667
rect 25421 24633 25455 24667
rect 31217 24633 31251 24667
rect 4537 24565 4571 24599
rect 7113 24565 7147 24599
rect 7297 24565 7331 24599
rect 13369 24565 13403 24599
rect 16037 24565 16071 24599
rect 19073 24565 19107 24599
rect 22109 24565 22143 24599
rect 22845 24565 22879 24599
rect 30113 24565 30147 24599
rect 7573 24361 7607 24395
rect 8217 24361 8251 24395
rect 8401 24361 8435 24395
rect 9137 24361 9171 24395
rect 10701 24361 10735 24395
rect 24777 24361 24811 24395
rect 26525 24361 26559 24395
rect 28365 24361 28399 24395
rect 32781 24361 32815 24395
rect 13553 24293 13587 24327
rect 6193 24225 6227 24259
rect 11897 24225 11931 24259
rect 21373 24225 21407 24259
rect 26065 24225 26099 24259
rect 3893 24157 3927 24191
rect 9781 24157 9815 24191
rect 12173 24157 12207 24191
rect 13185 24157 13219 24191
rect 15577 24157 15611 24191
rect 18705 24157 18739 24191
rect 19533 24157 19567 24191
rect 19625 24157 19659 24191
rect 19717 24157 19751 24191
rect 19901 24157 19935 24191
rect 20453 24157 20487 24191
rect 21931 24157 21965 24191
rect 23121 24157 23155 24191
rect 24409 24157 24443 24191
rect 25697 24157 25731 24191
rect 26801 24157 26835 24191
rect 26890 24154 26924 24188
rect 26985 24157 27019 24191
rect 27169 24157 27203 24191
rect 28365 24157 28399 24191
rect 28549 24157 28583 24191
rect 29561 24157 29595 24191
rect 31401 24157 31435 24191
rect 31657 24157 31691 24191
rect 4160 24089 4194 24123
rect 6460 24089 6494 24123
rect 8033 24089 8067 24123
rect 8953 24089 8987 24123
rect 10609 24089 10643 24123
rect 13369 24089 13403 24123
rect 17325 24089 17359 24123
rect 18521 24089 18555 24123
rect 20637 24089 20671 24123
rect 21189 24089 21223 24123
rect 22937 24089 22971 24123
rect 23673 24089 23707 24123
rect 24593 24089 24627 24123
rect 25881 24089 25915 24123
rect 29806 24089 29840 24123
rect 5273 24021 5307 24055
rect 8233 24021 8267 24055
rect 9153 24021 9187 24055
rect 9321 24021 9355 24055
rect 9965 24021 9999 24055
rect 19257 24021 19291 24055
rect 22109 24021 22143 24055
rect 23765 24021 23799 24055
rect 30941 24021 30975 24055
rect 5549 23817 5583 23851
rect 7757 23817 7791 23851
rect 9597 23817 9631 23851
rect 12081 23817 12115 23851
rect 25053 23817 25087 23851
rect 28273 23817 28307 23851
rect 29837 23817 29871 23851
rect 5181 23749 5215 23783
rect 5397 23749 5431 23783
rect 10425 23749 10459 23783
rect 10641 23749 10675 23783
rect 11713 23749 11747 23783
rect 14350 23749 14384 23783
rect 16957 23749 16991 23783
rect 19502 23749 19536 23783
rect 30757 23749 30791 23783
rect 4537 23681 4571 23715
rect 6377 23681 6411 23715
rect 6644 23681 6678 23715
rect 8217 23681 8251 23715
rect 8484 23681 8518 23715
rect 11897 23681 11931 23715
rect 13257 23681 13291 23715
rect 13350 23684 13384 23718
rect 13482 23681 13516 23715
rect 13645 23681 13679 23715
rect 14105 23681 14139 23715
rect 16773 23681 16807 23715
rect 17417 23681 17451 23715
rect 17673 23681 17707 23715
rect 19257 23681 19291 23715
rect 22109 23681 22143 23715
rect 23213 23681 23247 23715
rect 25329 23681 25363 23715
rect 25421 23681 25455 23715
rect 25513 23681 25547 23715
rect 25697 23681 25731 23715
rect 26157 23681 26191 23715
rect 26341 23681 26375 23715
rect 28529 23681 28563 23715
rect 28641 23681 28675 23715
rect 28733 23681 28767 23715
rect 28917 23681 28951 23715
rect 29469 23681 29503 23715
rect 29653 23681 29687 23715
rect 30389 23681 30423 23715
rect 30482 23681 30516 23715
rect 30665 23681 30699 23715
rect 30895 23681 30929 23715
rect 21833 23613 21867 23647
rect 15485 23545 15519 23579
rect 18797 23545 18831 23579
rect 20637 23545 20671 23579
rect 26157 23545 26191 23579
rect 4353 23477 4387 23511
rect 5365 23477 5399 23511
rect 10609 23477 10643 23511
rect 10793 23477 10827 23511
rect 13001 23477 13035 23511
rect 23305 23477 23339 23511
rect 31033 23477 31067 23511
rect 6745 23273 6779 23307
rect 8217 23273 8251 23307
rect 10701 23273 10735 23307
rect 11253 23273 11287 23307
rect 14657 23273 14691 23307
rect 17049 23273 17083 23307
rect 18613 23273 18647 23307
rect 21005 23273 21039 23307
rect 25605 23273 25639 23307
rect 26249 23273 26283 23307
rect 28457 23273 28491 23307
rect 9321 23137 9355 23171
rect 16313 23137 16347 23171
rect 3801 23069 3835 23103
rect 4068 23069 4102 23103
rect 6929 23069 6963 23103
rect 8401 23069 8435 23103
rect 11437 23069 11471 23103
rect 14289 23069 14323 23103
rect 16129 23069 16163 23103
rect 17279 23069 17313 23103
rect 17417 23069 17451 23103
rect 17509 23069 17543 23103
rect 17693 23069 17727 23103
rect 18429 23069 18463 23103
rect 19901 23069 19935 23103
rect 22109 23069 22143 23103
rect 22201 23069 22235 23103
rect 22293 23069 22327 23103
rect 22477 23069 22511 23103
rect 25237 23069 25271 23103
rect 25421 23069 25455 23103
rect 28089 23069 28123 23103
rect 28273 23069 28307 23103
rect 32689 23069 32723 23103
rect 9588 23001 9622 23035
rect 14473 23001 14507 23035
rect 15945 23001 15979 23035
rect 19717 23001 19751 23035
rect 20361 23001 20395 23035
rect 20913 23001 20947 23035
rect 26157 23001 26191 23035
rect 5181 22933 5215 22967
rect 20085 22933 20119 22967
rect 21833 22933 21867 22967
rect 32505 22933 32539 22967
rect 14381 22729 14415 22763
rect 20729 22729 20763 22763
rect 23213 22729 23247 22763
rect 23765 22729 23799 22763
rect 26433 22729 26467 22763
rect 4537 22661 4571 22695
rect 4753 22661 4787 22695
rect 6561 22661 6595 22695
rect 6777 22661 6811 22695
rect 11529 22661 11563 22695
rect 11729 22661 11763 22695
rect 19441 22661 19475 22695
rect 32404 22661 32438 22695
rect 7573 22593 7607 22627
rect 8309 22593 8343 22627
rect 10241 22593 10275 22627
rect 12541 22593 12575 22627
rect 13257 22593 13291 22627
rect 17509 22593 17543 22627
rect 18337 22593 18371 22627
rect 21833 22593 21867 22627
rect 22089 22593 22123 22627
rect 23673 22593 23707 22627
rect 23857 22593 23891 22627
rect 25053 22593 25087 22627
rect 25309 22593 25343 22627
rect 27721 22593 27755 22627
rect 27813 22593 27847 22627
rect 27905 22593 27939 22627
rect 28089 22593 28123 22627
rect 30205 22593 30239 22627
rect 30472 22593 30506 22627
rect 32137 22593 32171 22627
rect 34161 22593 34195 22627
rect 8585 22525 8619 22559
rect 13001 22525 13035 22559
rect 18153 22525 18187 22559
rect 4905 22457 4939 22491
rect 7389 22457 7423 22491
rect 10057 22457 10091 22491
rect 4721 22389 4755 22423
rect 6745 22389 6779 22423
rect 6929 22389 6963 22423
rect 11713 22389 11747 22423
rect 11897 22389 11931 22423
rect 12357 22389 12391 22423
rect 17601 22389 17635 22423
rect 18521 22389 18555 22423
rect 27445 22389 27479 22423
rect 31585 22389 31619 22423
rect 33517 22389 33551 22423
rect 33977 22389 34011 22423
rect 7021 22185 7055 22219
rect 12173 22185 12207 22219
rect 12817 22185 12851 22219
rect 18521 22185 18555 22219
rect 28825 22185 28859 22219
rect 30941 22185 30975 22219
rect 21189 22117 21223 22151
rect 7481 22049 7515 22083
rect 22477 22049 22511 22083
rect 29837 22049 29871 22083
rect 32965 22049 32999 22083
rect 34069 22049 34103 22083
rect 5641 21981 5675 22015
rect 7757 21981 7791 22015
rect 10793 21981 10827 22015
rect 14657 21981 14691 22015
rect 16497 21981 16531 22015
rect 19809 21981 19843 22015
rect 24593 21981 24627 22015
rect 24741 21981 24775 22015
rect 24961 21981 24995 22015
rect 25099 21981 25133 22015
rect 25697 21981 25731 22015
rect 25845 21981 25879 22015
rect 26065 21981 26099 22015
rect 26162 21981 26196 22015
rect 27445 21981 27479 22015
rect 30113 21981 30147 22015
rect 30205 21981 30239 22015
rect 30302 21981 30336 22015
rect 30481 21981 30515 22015
rect 31217 21981 31251 22015
rect 31309 21981 31343 22015
rect 31401 21981 31435 22015
rect 31585 21981 31619 22015
rect 32689 21981 32723 22015
rect 32873 21981 32907 22015
rect 33885 21981 33919 22015
rect 34161 21981 34195 22015
rect 5908 21913 5942 21947
rect 11060 21913 11094 21947
rect 12633 21913 12667 21947
rect 14924 21913 14958 21947
rect 16742 21913 16776 21947
rect 18337 21913 18371 21947
rect 20076 21913 20110 21947
rect 21833 21913 21867 21947
rect 22744 21913 22778 21947
rect 24869 21913 24903 21947
rect 25973 21913 26007 21947
rect 27701 21913 27735 21947
rect 12833 21845 12867 21879
rect 13001 21845 13035 21879
rect 16037 21845 16071 21879
rect 17877 21845 17911 21879
rect 18537 21845 18571 21879
rect 18705 21845 18739 21879
rect 21925 21845 21959 21879
rect 23857 21845 23891 21879
rect 25237 21845 25271 21879
rect 26341 21845 26375 21879
rect 32505 21845 32539 21879
rect 33701 21845 33735 21879
rect 7865 21641 7899 21675
rect 8493 21641 8527 21675
rect 12909 21641 12943 21675
rect 15577 21641 15611 21675
rect 18797 21641 18831 21675
rect 22293 21641 22327 21675
rect 22845 21641 22879 21675
rect 25329 21641 25363 21675
rect 27445 21641 27479 21675
rect 31033 21641 31067 21675
rect 32689 21641 32723 21675
rect 34989 21641 35023 21675
rect 7665 21573 7699 21607
rect 11796 21573 11830 21607
rect 15117 21573 15151 21607
rect 16773 21573 16807 21607
rect 21925 21573 21959 21607
rect 22141 21573 22175 21607
rect 28181 21573 28215 21607
rect 30205 21573 30239 21607
rect 32321 21573 32355 21607
rect 33876 21573 33910 21607
rect 4445 21505 4479 21539
rect 5089 21505 5123 21539
rect 6377 21505 6411 21539
rect 8677 21505 8711 21539
rect 9229 21505 9263 21539
rect 14933 21505 14967 21539
rect 15761 21505 15795 21539
rect 15853 21505 15887 21539
rect 16037 21505 16071 21539
rect 16129 21505 16163 21539
rect 17417 21505 17451 21539
rect 17684 21505 17718 21539
rect 19441 21505 19475 21539
rect 23121 21505 23155 21539
rect 23213 21505 23247 21539
rect 23305 21505 23339 21539
rect 23489 21505 23523 21539
rect 24041 21505 24075 21539
rect 27077 21505 27111 21539
rect 27261 21505 27295 21539
rect 27905 21505 27939 21539
rect 27998 21505 28032 21539
rect 28273 21505 28307 21539
rect 28370 21505 28404 21539
rect 29009 21505 29043 21539
rect 29193 21505 29227 21539
rect 29837 21505 29871 21539
rect 29985 21505 30019 21539
rect 30113 21505 30147 21539
rect 30343 21505 30377 21539
rect 30941 21505 30975 21539
rect 31125 21505 31159 21539
rect 32505 21505 32539 21539
rect 6653 21437 6687 21471
rect 11529 21437 11563 21471
rect 14749 21437 14783 21471
rect 16957 21437 16991 21471
rect 19717 21437 19751 21471
rect 29377 21437 29411 21471
rect 33609 21437 33643 21471
rect 4261 21301 4295 21335
rect 4905 21301 4939 21335
rect 7849 21301 7883 21335
rect 8033 21301 8067 21335
rect 10517 21301 10551 21335
rect 22109 21301 22143 21335
rect 28549 21301 28583 21335
rect 30481 21301 30515 21335
rect 6285 21097 6319 21131
rect 7573 21097 7607 21131
rect 7757 21097 7791 21131
rect 11345 21097 11379 21131
rect 12817 21097 12851 21131
rect 16221 21097 16255 21131
rect 18429 21097 18463 21131
rect 22661 21097 22695 21131
rect 23489 21097 23523 21131
rect 29929 21097 29963 21131
rect 31953 21097 31987 21131
rect 33977 21097 34011 21131
rect 26525 21029 26559 21063
rect 27261 21029 27295 21063
rect 8953 20961 8987 20995
rect 14105 20961 14139 20995
rect 21005 20961 21039 20995
rect 3801 20893 3835 20927
rect 4068 20893 4102 20927
rect 6469 20893 6503 20927
rect 8401 20893 8435 20927
rect 11529 20893 11563 20927
rect 12725 20893 12759 20927
rect 16405 20893 16439 20927
rect 16497 20893 16531 20927
rect 16681 20893 16715 20927
rect 16773 20893 16807 20927
rect 17785 20893 17819 20927
rect 19257 20893 19291 20927
rect 19533 20893 19567 20927
rect 21281 20893 21315 20927
rect 22293 20893 22327 20927
rect 23121 20893 23155 20927
rect 24409 20893 24443 20927
rect 24502 20893 24536 20927
rect 24777 20893 24811 20927
rect 24915 20893 24949 20927
rect 27813 20893 27847 20927
rect 29561 20893 29595 20927
rect 29745 20893 29779 20927
rect 30573 20893 30607 20927
rect 30829 20893 30863 20927
rect 7389 20825 7423 20859
rect 9220 20825 9254 20859
rect 14372 20825 14406 20859
rect 22477 20825 22511 20859
rect 23305 20825 23339 20859
rect 24685 20825 24719 20859
rect 25605 20825 25639 20859
rect 26341 20825 26375 20859
rect 27077 20825 27111 20859
rect 27997 20825 28031 20859
rect 33609 20825 33643 20859
rect 33793 20825 33827 20859
rect 5181 20757 5215 20791
rect 7589 20757 7623 20791
rect 8217 20757 8251 20791
rect 10333 20757 10367 20791
rect 15485 20757 15519 20791
rect 25053 20757 25087 20791
rect 25697 20757 25731 20791
rect 28181 20757 28215 20791
rect 5565 20553 5599 20587
rect 5733 20553 5767 20587
rect 6577 20553 6611 20587
rect 6745 20553 6779 20587
rect 10425 20553 10459 20587
rect 11713 20553 11747 20587
rect 14749 20553 14783 20587
rect 17693 20553 17727 20587
rect 19809 20553 19843 20587
rect 24593 20553 24627 20587
rect 27905 20553 27939 20587
rect 28457 20553 28491 20587
rect 3792 20485 3826 20519
rect 5365 20485 5399 20519
rect 6377 20485 6411 20519
rect 7389 20485 7423 20519
rect 7589 20485 7623 20519
rect 14105 20485 14139 20519
rect 16865 20485 16899 20519
rect 18889 20485 18923 20519
rect 25513 20485 25547 20519
rect 26985 20485 27019 20519
rect 29828 20485 29862 20519
rect 3065 20417 3099 20451
rect 8585 20417 8619 20451
rect 8841 20417 8875 20451
rect 10609 20417 10643 20451
rect 11529 20417 11563 20451
rect 13369 20417 13403 20451
rect 14933 20417 14967 20451
rect 15025 20417 15059 20451
rect 15209 20417 15243 20451
rect 15301 20417 15335 20451
rect 15853 20417 15887 20451
rect 15945 20417 15979 20451
rect 16681 20417 16715 20451
rect 17877 20417 17911 20451
rect 17969 20417 18003 20451
rect 18153 20417 18187 20451
rect 18245 20417 18279 20451
rect 18705 20417 18739 20451
rect 20085 20417 20119 20451
rect 20177 20417 20211 20451
rect 20269 20417 20303 20451
rect 20453 20417 20487 20451
rect 22661 20417 22695 20451
rect 22845 20417 22879 20451
rect 24501 20417 24535 20451
rect 24685 20417 24719 20451
rect 25145 20417 25179 20451
rect 25238 20417 25272 20451
rect 25421 20417 25455 20451
rect 25651 20417 25685 20451
rect 27169 20417 27203 20451
rect 27813 20417 27847 20451
rect 27997 20417 28031 20451
rect 28733 20417 28767 20451
rect 28825 20417 28859 20451
rect 28917 20417 28951 20451
rect 29101 20417 29135 20451
rect 32505 20417 32539 20451
rect 33977 20417 34011 20451
rect 34897 20417 34931 20451
rect 3525 20349 3559 20383
rect 14289 20349 14323 20383
rect 29561 20349 29595 20383
rect 32781 20349 32815 20383
rect 34253 20349 34287 20383
rect 13461 20281 13495 20315
rect 32689 20281 32723 20315
rect 34161 20281 34195 20315
rect 2881 20213 2915 20247
rect 4905 20213 4939 20247
rect 5549 20213 5583 20247
rect 6561 20213 6595 20247
rect 7573 20213 7607 20247
rect 7757 20213 7791 20247
rect 9965 20213 9999 20247
rect 16129 20213 16163 20247
rect 17049 20213 17083 20247
rect 19073 20213 19107 20247
rect 23029 20213 23063 20247
rect 25789 20213 25823 20247
rect 27353 20213 27387 20247
rect 30941 20213 30975 20247
rect 32321 20213 32355 20247
rect 33793 20213 33827 20247
rect 34713 20213 34747 20247
rect 5181 20009 5215 20043
rect 7573 20009 7607 20043
rect 8217 20009 8251 20043
rect 10333 20009 10367 20043
rect 31401 20009 31435 20043
rect 33701 20009 33735 20043
rect 7757 19941 7791 19975
rect 8953 19873 8987 19907
rect 19901 19873 19935 19907
rect 21741 19873 21775 19907
rect 22017 19873 22051 19907
rect 32321 19873 32355 19907
rect 3801 19805 3835 19839
rect 4057 19805 4091 19839
rect 6929 19805 6963 19839
rect 8401 19805 8435 19839
rect 9209 19805 9243 19839
rect 10977 19805 11011 19839
rect 15485 19805 15519 19839
rect 15577 19805 15611 19839
rect 15669 19805 15703 19839
rect 15853 19805 15887 19839
rect 16865 19805 16899 19839
rect 18245 19805 18279 19839
rect 18334 19805 18368 19839
rect 18429 19805 18463 19839
rect 18613 19805 18647 19839
rect 23305 19805 23339 19839
rect 23397 19805 23431 19839
rect 23489 19805 23523 19839
rect 23673 19805 23707 19839
rect 24409 19805 24443 19839
rect 24502 19805 24536 19839
rect 24874 19805 24908 19839
rect 26341 19805 26375 19839
rect 26489 19805 26523 19839
rect 26709 19805 26743 19839
rect 26847 19805 26881 19839
rect 27701 19805 27735 19839
rect 27813 19805 27847 19839
rect 27905 19805 27939 19839
rect 28089 19805 28123 19839
rect 30113 19805 30147 19839
rect 34713 19805 34747 19839
rect 34897 19805 34931 19839
rect 7389 19737 7423 19771
rect 7589 19737 7623 19771
rect 11222 19737 11256 19771
rect 14105 19737 14139 19771
rect 14289 19737 14323 19771
rect 16681 19737 16715 19771
rect 20168 19737 20202 19771
rect 24685 19737 24719 19771
rect 24777 19737 24811 19771
rect 26617 19737 26651 19771
rect 32566 19737 32600 19771
rect 6745 19669 6779 19703
rect 12357 19669 12391 19703
rect 14473 19669 14507 19703
rect 15209 19669 15243 19703
rect 17049 19669 17083 19703
rect 17969 19669 18003 19703
rect 21281 19669 21315 19703
rect 23029 19669 23063 19703
rect 25053 19669 25087 19703
rect 26985 19669 27019 19703
rect 27445 19669 27479 19703
rect 35081 19669 35115 19703
rect 4997 19465 5031 19499
rect 5641 19465 5675 19499
rect 9965 19465 9999 19499
rect 13185 19465 13219 19499
rect 15485 19465 15519 19499
rect 18705 19465 18739 19499
rect 20453 19465 20487 19499
rect 28365 19465 28399 19499
rect 30205 19465 30239 19499
rect 32229 19465 32263 19499
rect 33333 19465 33367 19499
rect 35173 19465 35207 19499
rect 4629 19397 4663 19431
rect 4845 19397 4879 19431
rect 6622 19397 6656 19431
rect 11897 19397 11931 19431
rect 14372 19397 14406 19431
rect 19165 19397 19199 19431
rect 22560 19397 22594 19431
rect 29070 19397 29104 19431
rect 5825 19329 5859 19363
rect 6377 19329 6411 19363
rect 8585 19329 8619 19363
rect 8841 19329 8875 19363
rect 10609 19329 10643 19363
rect 10793 19329 10827 19363
rect 14105 19329 14139 19363
rect 15945 19329 15979 19363
rect 16129 19329 16163 19363
rect 16681 19329 16715 19363
rect 16865 19329 16899 19363
rect 17325 19329 17359 19363
rect 17592 19329 17626 19363
rect 22293 19329 22327 19363
rect 24133 19329 24167 19363
rect 24400 19329 24434 19363
rect 26985 19329 27019 19363
rect 27241 19329 27275 19363
rect 28825 19329 28859 19363
rect 30941 19329 30975 19363
rect 32413 19329 32447 19363
rect 33149 19329 33183 19363
rect 33793 19329 33827 19363
rect 34060 19329 34094 19363
rect 37565 19329 37599 19363
rect 32965 19261 32999 19295
rect 37289 19261 37323 19295
rect 16681 19193 16715 19227
rect 23673 19193 23707 19227
rect 4813 19125 4847 19159
rect 7757 19125 7791 19159
rect 10977 19125 11011 19159
rect 16037 19125 16071 19159
rect 25513 19125 25547 19159
rect 30757 19125 30791 19159
rect 5457 18921 5491 18955
rect 6653 18921 6687 18955
rect 8125 18921 8159 18955
rect 10333 18921 10367 18955
rect 23213 18921 23247 18955
rect 24409 18921 24443 18955
rect 26525 18921 26559 18955
rect 27997 18921 28031 18955
rect 34069 18921 34103 18955
rect 6837 18853 6871 18887
rect 14381 18785 14415 18819
rect 19809 18785 19843 18819
rect 22569 18785 22603 18819
rect 32597 18785 32631 18819
rect 34713 18785 34747 18819
rect 4169 18717 4203 18751
rect 8309 18717 8343 18751
rect 10609 18717 10643 18751
rect 10701 18717 10735 18751
rect 10793 18717 10827 18751
rect 10977 18717 11011 18751
rect 11713 18717 11747 18751
rect 11805 18717 11839 18751
rect 11897 18717 11931 18751
rect 12081 18717 12115 18751
rect 13185 18717 13219 18751
rect 13277 18717 13311 18751
rect 13369 18717 13403 18751
rect 13553 18717 13587 18751
rect 14105 18717 14139 18751
rect 15761 18717 15795 18751
rect 15853 18717 15887 18751
rect 15945 18717 15979 18751
rect 16129 18717 16163 18751
rect 16865 18717 16899 18751
rect 16957 18717 16991 18751
rect 17049 18717 17083 18751
rect 17233 18717 17267 18751
rect 18337 18717 18371 18751
rect 18429 18717 18463 18751
rect 18521 18717 18555 18751
rect 18705 18717 18739 18751
rect 20085 18717 20119 18751
rect 21327 18717 21361 18751
rect 21446 18714 21480 18748
rect 21557 18717 21591 18751
rect 21753 18717 21787 18751
rect 22385 18717 22419 18751
rect 24685 18717 24719 18751
rect 24777 18717 24811 18751
rect 24869 18717 24903 18751
rect 25053 18717 25087 18751
rect 26801 18717 26835 18751
rect 26893 18717 26927 18751
rect 26985 18717 27019 18751
rect 27169 18717 27203 18751
rect 27629 18717 27663 18751
rect 27813 18717 27847 18751
rect 30665 18717 30699 18751
rect 30921 18717 30955 18751
rect 32781 18717 32815 18751
rect 33885 18717 33919 18751
rect 34989 18717 35023 18751
rect 6469 18649 6503 18683
rect 22201 18649 22235 18683
rect 23121 18649 23155 18683
rect 33701 18649 33735 18683
rect 6669 18581 6703 18615
rect 11437 18581 11471 18615
rect 12909 18581 12943 18615
rect 15485 18581 15519 18615
rect 16589 18581 16623 18615
rect 18061 18581 18095 18615
rect 21097 18581 21131 18615
rect 32045 18581 32079 18615
rect 32965 18581 32999 18615
rect 7941 18377 7975 18411
rect 10977 18377 11011 18411
rect 12081 18377 12115 18411
rect 18153 18377 18187 18411
rect 19901 18377 19935 18411
rect 32505 18377 32539 18411
rect 11897 18309 11931 18343
rect 21097 18309 21131 18343
rect 21281 18309 21315 18343
rect 23121 18309 23155 18343
rect 24317 18309 24351 18343
rect 25145 18309 25179 18343
rect 32321 18309 32355 18343
rect 7849 18241 7883 18275
rect 9597 18241 9631 18275
rect 9864 18241 9898 18275
rect 11713 18241 11747 18275
rect 12633 18241 12667 18275
rect 14611 18241 14645 18275
rect 14749 18241 14783 18275
rect 14862 18244 14896 18278
rect 15025 18241 15059 18275
rect 15577 18241 15611 18275
rect 17417 18241 17451 18275
rect 17601 18241 17635 18275
rect 18383 18241 18417 18275
rect 18521 18241 18555 18275
rect 18613 18241 18647 18275
rect 18797 18241 18831 18275
rect 20177 18241 20211 18275
rect 20269 18241 20303 18275
rect 20361 18241 20395 18275
rect 20545 18241 20579 18275
rect 21833 18241 21867 18275
rect 22017 18241 22051 18275
rect 23305 18241 23339 18275
rect 24133 18241 24167 18275
rect 30665 18241 30699 18275
rect 30941 18241 30975 18275
rect 32137 18241 32171 18275
rect 33057 18241 33091 18275
rect 33333 18173 33367 18207
rect 37289 18173 37323 18207
rect 37565 18173 37599 18207
rect 12817 18105 12851 18139
rect 22201 18105 22235 18139
rect 24501 18105 24535 18139
rect 14381 18037 14415 18071
rect 15669 18037 15703 18071
rect 25237 18037 25271 18071
rect 30481 18037 30515 18071
rect 30849 18037 30883 18071
rect 9505 17833 9539 17867
rect 11805 17833 11839 17867
rect 15853 17833 15887 17867
rect 19625 17833 19659 17867
rect 22569 17833 22603 17867
rect 30849 17833 30883 17867
rect 33425 17833 33459 17867
rect 6929 17765 6963 17799
rect 15209 17765 15243 17799
rect 12909 17697 12943 17731
rect 21189 17697 21223 17731
rect 23029 17697 23063 17731
rect 24869 17697 24903 17731
rect 28457 17697 28491 17731
rect 28641 17697 28675 17731
rect 31585 17697 31619 17731
rect 6469 17629 6503 17663
rect 7113 17629 7147 17663
rect 10977 17629 11011 17663
rect 11069 17629 11103 17663
rect 11161 17629 11195 17663
rect 11345 17629 11379 17663
rect 12081 17629 12115 17663
rect 12173 17629 12207 17663
rect 12265 17629 12299 17663
rect 12449 17629 12483 17663
rect 13093 17629 13127 17663
rect 16497 17629 16531 17663
rect 19441 17629 19475 17663
rect 20361 17629 20395 17663
rect 20453 17629 20487 17663
rect 20545 17629 20579 17663
rect 20729 17629 20763 17663
rect 23213 17629 23247 17663
rect 28365 17629 28399 17663
rect 29653 17629 29687 17663
rect 30481 17629 30515 17663
rect 31861 17629 31895 17663
rect 33057 17629 33091 17663
rect 33241 17629 33275 17663
rect 34713 17629 34747 17663
rect 9413 17561 9447 17595
rect 15025 17561 15059 17595
rect 15761 17561 15795 17595
rect 17233 17561 17267 17595
rect 19257 17561 19291 17595
rect 21456 17561 21490 17595
rect 25136 17561 25170 17595
rect 29837 17561 29871 17595
rect 30665 17561 30699 17595
rect 34958 17561 34992 17595
rect 6285 17493 6319 17527
rect 10701 17493 10735 17527
rect 13277 17493 13311 17527
rect 16589 17493 16623 17527
rect 17325 17493 17359 17527
rect 20085 17493 20119 17527
rect 23397 17493 23431 17527
rect 26249 17493 26283 17527
rect 28641 17493 28675 17527
rect 30021 17493 30055 17527
rect 36093 17493 36127 17527
rect 7205 17289 7239 17323
rect 12541 17289 12575 17323
rect 13461 17289 13495 17323
rect 18383 17289 18417 17323
rect 22569 17289 22603 17323
rect 26985 17289 27019 17323
rect 29285 17289 29319 17323
rect 6561 17221 6595 17255
rect 6745 17221 6779 17255
rect 11713 17221 11747 17255
rect 13185 17221 13219 17255
rect 14381 17221 14415 17255
rect 24961 17221 24995 17255
rect 32321 17221 32355 17255
rect 34958 17221 34992 17255
rect 2964 17153 2998 17187
rect 5825 17153 5859 17187
rect 6377 17153 6411 17187
rect 7389 17153 7423 17187
rect 8033 17153 8067 17187
rect 8677 17153 8711 17187
rect 12357 17153 12391 17187
rect 14105 17153 14139 17187
rect 14197 17153 14231 17187
rect 15117 17153 15151 17187
rect 15209 17153 15243 17187
rect 15393 17153 15427 17187
rect 15485 17153 15519 17187
rect 15945 17153 15979 17187
rect 17141 17153 17175 17187
rect 17325 17153 17359 17187
rect 19717 17153 19751 17187
rect 19809 17153 19843 17187
rect 19901 17153 19935 17187
rect 20079 17153 20113 17187
rect 20821 17153 20855 17187
rect 20913 17153 20947 17187
rect 21005 17153 21039 17187
rect 21189 17153 21223 17187
rect 21925 17153 21959 17187
rect 23305 17153 23339 17187
rect 23581 17153 23615 17187
rect 24593 17153 24627 17187
rect 24777 17153 24811 17187
rect 25881 17153 25915 17187
rect 26157 17153 26191 17187
rect 27169 17153 27203 17187
rect 28172 17153 28206 17187
rect 29745 17153 29779 17187
rect 30001 17153 30035 17187
rect 32137 17153 32171 17187
rect 33149 17153 33183 17187
rect 33793 17153 33827 17187
rect 2697 17085 2731 17119
rect 18153 17085 18187 17119
rect 19441 17085 19475 17119
rect 27905 17085 27939 17119
rect 34713 17085 34747 17119
rect 5641 17017 5675 17051
rect 7849 17017 7883 17051
rect 11897 17017 11931 17051
rect 26065 17017 26099 17051
rect 32965 17017 32999 17051
rect 4077 16949 4111 16983
rect 8493 16949 8527 16983
rect 14933 16949 14967 16983
rect 16037 16949 16071 16983
rect 17233 16949 17267 16983
rect 20545 16949 20579 16983
rect 25697 16949 25731 16983
rect 31125 16949 31159 16983
rect 32505 16949 32539 16983
rect 33609 16949 33643 16983
rect 36093 16949 36127 16983
rect 7389 16745 7423 16779
rect 9321 16745 9355 16779
rect 24777 16745 24811 16779
rect 29745 16745 29779 16779
rect 5181 16677 5215 16711
rect 21465 16677 21499 16711
rect 31677 16677 31711 16711
rect 33793 16677 33827 16711
rect 3801 16609 3835 16643
rect 6561 16609 6595 16643
rect 19257 16609 19291 16643
rect 22477 16609 22511 16643
rect 24869 16609 24903 16643
rect 26065 16609 26099 16643
rect 27261 16609 27295 16643
rect 30389 16609 30423 16643
rect 30849 16609 30883 16643
rect 32505 16609 32539 16643
rect 33333 16609 33367 16643
rect 1869 16541 1903 16575
rect 4068 16541 4102 16575
rect 7205 16541 7239 16575
rect 8217 16541 8251 16575
rect 8401 16541 8435 16575
rect 11023 16541 11057 16575
rect 11158 16541 11192 16575
rect 11258 16541 11292 16575
rect 11437 16541 11471 16575
rect 13185 16541 13219 16575
rect 13274 16538 13308 16572
rect 13369 16541 13403 16575
rect 13565 16541 13599 16575
rect 14933 16541 14967 16575
rect 15025 16541 15059 16575
rect 15117 16541 15151 16575
rect 15301 16541 15335 16575
rect 15761 16541 15795 16575
rect 16865 16541 16899 16575
rect 16957 16541 16991 16575
rect 17054 16541 17088 16575
rect 17233 16541 17267 16575
rect 17877 16541 17911 16575
rect 17969 16541 18003 16575
rect 18153 16541 18187 16575
rect 18245 16541 18279 16575
rect 19524 16541 19558 16575
rect 21649 16541 21683 16575
rect 21741 16541 21775 16575
rect 21925 16541 21959 16575
rect 22017 16541 22051 16575
rect 24593 16541 24627 16575
rect 25881 16541 25915 16575
rect 29929 16541 29963 16575
rect 30573 16541 30607 16575
rect 30757 16541 30791 16575
rect 31309 16541 31343 16575
rect 32321 16541 32355 16575
rect 33977 16541 34011 16575
rect 2136 16473 2170 16507
rect 6193 16473 6227 16507
rect 6377 16473 6411 16507
rect 7021 16473 7055 16507
rect 8309 16473 8343 16507
rect 8953 16473 8987 16507
rect 9137 16473 9171 16507
rect 22744 16473 22778 16507
rect 27528 16473 27562 16507
rect 31493 16473 31527 16507
rect 32137 16473 32171 16507
rect 32965 16473 32999 16507
rect 33149 16473 33183 16507
rect 35081 16473 35115 16507
rect 3249 16405 3283 16439
rect 10793 16405 10827 16439
rect 12909 16405 12943 16439
rect 14657 16405 14691 16439
rect 15945 16405 15979 16439
rect 16589 16405 16623 16439
rect 17693 16405 17727 16439
rect 20637 16405 20671 16439
rect 23857 16405 23891 16439
rect 24409 16405 24443 16439
rect 28641 16405 28675 16439
rect 36369 16405 36403 16439
rect 4077 16201 4111 16235
rect 6745 16201 6779 16235
rect 9321 16201 9355 16235
rect 15669 16201 15703 16235
rect 19993 16201 20027 16235
rect 22017 16201 22051 16235
rect 28825 16201 28859 16235
rect 34069 16201 34103 16235
rect 36369 16201 36403 16235
rect 5641 16133 5675 16167
rect 5825 16133 5859 16167
rect 6561 16133 6595 16167
rect 8208 16133 8242 16167
rect 14556 16133 14590 16167
rect 18705 16133 18739 16167
rect 19625 16133 19659 16167
rect 19809 16133 19843 16167
rect 21925 16133 21959 16167
rect 23213 16133 23247 16167
rect 23397 16133 23431 16167
rect 27537 16133 27571 16167
rect 31217 16133 31251 16167
rect 31401 16133 31435 16167
rect 32956 16133 32990 16167
rect 2697 16065 2731 16099
rect 2964 16065 2998 16099
rect 4997 16065 5031 16099
rect 5457 16065 5491 16099
rect 6377 16065 6411 16099
rect 7389 16065 7423 16099
rect 10609 16065 10643 16099
rect 10698 16065 10732 16099
rect 10798 16065 10832 16099
rect 10977 16065 11011 16099
rect 12440 16065 12474 16099
rect 16773 16065 16807 16099
rect 17040 16065 17074 16099
rect 18613 16065 18647 16099
rect 20637 16065 20671 16099
rect 20821 16065 20855 16099
rect 22569 16065 22603 16099
rect 22753 16065 22787 16099
rect 24133 16065 24167 16099
rect 25320 16065 25354 16099
rect 27169 16065 27203 16099
rect 27997 16065 28031 16099
rect 28733 16065 28767 16099
rect 28917 16065 28951 16099
rect 30389 16065 30423 16099
rect 30573 16065 30607 16099
rect 34529 16065 34563 16099
rect 34785 16065 34819 16099
rect 36553 16065 36587 16099
rect 7941 15997 7975 16031
rect 12173 15997 12207 16031
rect 14289 15997 14323 16031
rect 25053 15997 25087 16031
rect 26985 15997 27019 16031
rect 28089 15997 28123 16031
rect 28273 15997 28307 16031
rect 32689 15997 32723 16031
rect 18153 15929 18187 15963
rect 24317 15929 24351 15963
rect 26433 15929 26467 15963
rect 4813 15861 4847 15895
rect 7205 15861 7239 15895
rect 10333 15861 10367 15895
rect 13553 15861 13587 15895
rect 20729 15861 20763 15895
rect 22569 15861 22603 15895
rect 23581 15861 23615 15895
rect 27445 15861 27479 15895
rect 28181 15861 28215 15895
rect 30757 15861 30791 15895
rect 31585 15861 31619 15895
rect 35909 15861 35943 15895
rect 3249 15657 3283 15691
rect 12725 15657 12759 15691
rect 14933 15657 14967 15691
rect 15485 15657 15519 15691
rect 17693 15657 17727 15691
rect 19809 15657 19843 15691
rect 23305 15657 23339 15691
rect 26157 15657 26191 15691
rect 27629 15657 27663 15691
rect 36093 15657 36127 15691
rect 11989 15589 12023 15623
rect 31493 15589 31527 15623
rect 34161 15589 34195 15623
rect 1869 15521 1903 15555
rect 36553 15521 36587 15555
rect 3801 15453 3835 15487
rect 5641 15453 5675 15487
rect 7665 15453 7699 15487
rect 9137 15453 9171 15487
rect 9781 15453 9815 15487
rect 10048 15453 10082 15487
rect 13001 15453 13035 15487
rect 13093 15453 13127 15487
rect 13185 15453 13219 15487
rect 13369 15453 13403 15487
rect 14841 15453 14875 15487
rect 15025 15453 15059 15487
rect 15485 15453 15519 15487
rect 15669 15453 15703 15487
rect 17693 15453 17727 15487
rect 17877 15453 17911 15487
rect 20913 15453 20947 15487
rect 21005 15453 21039 15487
rect 21097 15453 21131 15487
rect 21281 15453 21315 15487
rect 21925 15453 21959 15487
rect 22017 15453 22051 15487
rect 22201 15453 22235 15487
rect 22293 15453 22327 15487
rect 23489 15453 23523 15487
rect 24869 15453 24903 15487
rect 26157 15453 26191 15487
rect 26341 15453 26375 15487
rect 27629 15453 27663 15487
rect 27813 15453 27847 15487
rect 29837 15453 29871 15487
rect 30297 15453 30331 15487
rect 30481 15453 30515 15487
rect 30665 15453 30699 15487
rect 32137 15453 32171 15487
rect 32781 15453 32815 15487
rect 33048 15453 33082 15487
rect 34713 15453 34747 15487
rect 2136 15385 2170 15419
rect 4068 15385 4102 15419
rect 5908 15385 5942 15419
rect 7481 15385 7515 15419
rect 11621 15385 11655 15419
rect 11805 15385 11839 15419
rect 19717 15385 19751 15419
rect 31125 15385 31159 15419
rect 31309 15385 31343 15419
rect 31953 15385 31987 15419
rect 34958 15385 34992 15419
rect 36798 15385 36832 15419
rect 5181 15317 5215 15351
rect 7021 15317 7055 15351
rect 7849 15317 7883 15351
rect 8953 15317 8987 15351
rect 11161 15317 11195 15351
rect 20637 15317 20671 15351
rect 21741 15317 21775 15351
rect 24961 15317 24995 15351
rect 29653 15317 29687 15351
rect 32321 15317 32355 15351
rect 37933 15317 37967 15351
rect 4813 15113 4847 15147
rect 6745 15113 6779 15147
rect 8033 15113 8067 15147
rect 13369 15113 13403 15147
rect 17601 15113 17635 15147
rect 34069 15113 34103 15147
rect 36369 15113 36403 15147
rect 2964 15045 2998 15079
rect 7205 15045 7239 15079
rect 13001 15045 13035 15079
rect 13185 15045 13219 15079
rect 15209 15045 15243 15079
rect 16957 15045 16991 15079
rect 18521 15045 18555 15079
rect 32956 15045 32990 15079
rect 34785 15045 34819 15079
rect 2697 14977 2731 15011
rect 4997 14977 5031 15011
rect 5457 14977 5491 15011
rect 5641 14977 5675 15011
rect 6377 14977 6411 15011
rect 6561 14977 6595 15011
rect 7389 14977 7423 15011
rect 8217 14977 8251 15011
rect 8861 14977 8895 15011
rect 9505 14977 9539 15011
rect 10149 14977 10183 15011
rect 15945 14977 15979 15011
rect 18245 14977 18279 15011
rect 18337 14977 18371 15011
rect 19993 14977 20027 15011
rect 21833 14977 21867 15011
rect 22100 14977 22134 15011
rect 23673 14977 23707 15011
rect 23857 14977 23891 15011
rect 24041 14977 24075 15011
rect 24685 14977 24719 15011
rect 25605 14977 25639 15011
rect 28641 14977 28675 15011
rect 28825 14977 28859 15011
rect 30021 14977 30055 15011
rect 30849 14977 30883 15011
rect 34529 14977 34563 15011
rect 36553 14977 36587 15011
rect 15577 14909 15611 14943
rect 17325 14909 17359 14943
rect 19717 14909 19751 14943
rect 25421 14909 25455 14943
rect 29837 14909 29871 14943
rect 30665 14909 30699 14943
rect 32689 14909 32723 14943
rect 4077 14841 4111 14875
rect 9321 14841 9355 14875
rect 9965 14841 9999 14875
rect 5825 14773 5859 14807
rect 7573 14773 7607 14807
rect 8677 14773 8711 14807
rect 15347 14773 15381 14807
rect 15485 14773 15519 14807
rect 17095 14773 17129 14807
rect 17233 14773 17267 14807
rect 23213 14773 23247 14807
rect 24501 14773 24535 14807
rect 25789 14773 25823 14807
rect 28641 14773 28675 14807
rect 30205 14773 30239 14807
rect 31033 14773 31067 14807
rect 35909 14773 35943 14807
rect 3249 14569 3283 14603
rect 8217 14569 8251 14603
rect 13461 14569 13495 14603
rect 22017 14569 22051 14603
rect 26065 14569 26099 14603
rect 28089 14569 28123 14603
rect 28825 14569 28859 14603
rect 33793 14569 33827 14603
rect 16313 14501 16347 14535
rect 28917 14501 28951 14535
rect 3801 14433 3835 14467
rect 9781 14433 9815 14467
rect 28273 14433 28307 14467
rect 29009 14433 29043 14467
rect 29561 14433 29595 14467
rect 34713 14433 34747 14467
rect 1869 14365 1903 14399
rect 4068 14365 4102 14399
rect 5641 14365 5675 14399
rect 9137 14365 9171 14399
rect 12081 14365 12115 14399
rect 15117 14365 15151 14399
rect 15393 14365 15427 14399
rect 15761 14365 15795 14399
rect 16313 14365 16347 14399
rect 17509 14365 17543 14399
rect 17877 14365 17911 14399
rect 18061 14365 18095 14399
rect 18337 14365 18371 14399
rect 19257 14365 19291 14399
rect 19533 14365 19567 14399
rect 19993 14365 20027 14399
rect 20177 14365 20211 14399
rect 21925 14365 21959 14399
rect 23213 14365 23247 14399
rect 26985 14365 27019 14399
rect 27169 14365 27203 14399
rect 27997 14365 28031 14399
rect 28733 14365 28767 14399
rect 29817 14365 29851 14399
rect 31585 14365 31619 14399
rect 32321 14365 32355 14399
rect 32505 14365 32539 14399
rect 33977 14365 34011 14399
rect 34969 14365 35003 14399
rect 2136 14297 2170 14331
rect 7849 14297 7883 14331
rect 8033 14297 8067 14331
rect 10048 14297 10082 14331
rect 12348 14297 12382 14331
rect 19441 14297 19475 14331
rect 24777 14297 24811 14331
rect 32137 14297 32171 14331
rect 32965 14297 32999 14331
rect 33149 14297 33183 14331
rect 5181 14229 5215 14263
rect 6929 14229 6963 14263
rect 8953 14229 8987 14263
rect 11161 14229 11195 14263
rect 19355 14229 19389 14263
rect 20085 14229 20119 14263
rect 23397 14229 23431 14263
rect 27077 14229 27111 14263
rect 28273 14229 28307 14263
rect 30941 14229 30975 14263
rect 31401 14229 31435 14263
rect 33333 14229 33367 14263
rect 36093 14229 36127 14263
rect 4077 14025 4111 14059
rect 6745 14025 6779 14059
rect 7573 14025 7607 14059
rect 11621 14025 11655 14059
rect 13185 14025 13219 14059
rect 14197 14025 14231 14059
rect 16037 14025 16071 14059
rect 20453 14025 20487 14059
rect 29745 14025 29779 14059
rect 31401 14025 31435 14059
rect 32965 14025 32999 14059
rect 35909 14025 35943 14059
rect 2964 13957 2998 13991
rect 7389 13957 7423 13991
rect 9413 13957 9447 13991
rect 10149 13957 10183 13991
rect 12335 13957 12369 13991
rect 19340 13957 19374 13991
rect 32505 13957 32539 13991
rect 2697 13889 2731 13923
rect 5825 13889 5859 13923
rect 6377 13889 6411 13923
rect 6561 13889 6595 13923
rect 7205 13889 7239 13923
rect 8217 13889 8251 13923
rect 8401 13889 8435 13923
rect 9045 13889 9079 13923
rect 9229 13889 9263 13923
rect 10517 13889 10551 13923
rect 11529 13889 11563 13923
rect 11713 13889 11747 13923
rect 12633 13889 12667 13923
rect 13093 13889 13127 13923
rect 13277 13889 13311 13923
rect 13829 13889 13863 13923
rect 14933 13889 14967 13923
rect 15117 13889 15151 13923
rect 15485 13889 15519 13923
rect 15853 13889 15887 13923
rect 17141 13889 17175 13923
rect 17969 13889 18003 13923
rect 19073 13889 19107 13923
rect 21925 13889 21959 13923
rect 22109 13889 22143 13923
rect 22845 13889 22879 13923
rect 23112 13889 23146 13923
rect 24777 13889 24811 13923
rect 25044 13889 25078 13923
rect 27169 13889 27203 13923
rect 27436 13889 27470 13923
rect 29101 13889 29135 13923
rect 29929 13889 29963 13923
rect 31585 13889 31619 13923
rect 32137 13889 32171 13923
rect 32321 13889 32355 13923
rect 33149 13889 33183 13923
rect 33793 13889 33827 13923
rect 34529 13889 34563 13923
rect 34785 13889 34819 13923
rect 8585 13821 8619 13855
rect 10333 13821 10367 13855
rect 12449 13821 12483 13855
rect 13921 13821 13955 13855
rect 17877 13821 17911 13855
rect 5641 13753 5675 13787
rect 12265 13753 12299 13787
rect 17969 13753 18003 13787
rect 28549 13753 28583 13787
rect 33609 13753 33643 13787
rect 10333 13685 10367 13719
rect 10425 13685 10459 13719
rect 12541 13685 12575 13719
rect 14013 13685 14047 13719
rect 22017 13685 22051 13719
rect 24225 13685 24259 13719
rect 26157 13685 26191 13719
rect 29193 13685 29227 13719
rect 6285 13481 6319 13515
rect 9321 13481 9355 13515
rect 14197 13481 14231 13515
rect 17601 13481 17635 13515
rect 23673 13481 23707 13515
rect 24501 13481 24535 13515
rect 26433 13481 26467 13515
rect 27721 13481 27755 13515
rect 30941 13481 30975 13515
rect 33425 13481 33459 13515
rect 8401 13413 8435 13447
rect 13461 13413 13495 13447
rect 17233 13413 17267 13447
rect 18337 13413 18371 13447
rect 32781 13413 32815 13447
rect 12081 13345 12115 13379
rect 17325 13345 17359 13379
rect 19257 13345 19291 13379
rect 19717 13345 19751 13379
rect 24685 13345 24719 13379
rect 26341 13345 26375 13379
rect 26525 13345 26559 13379
rect 27077 13345 27111 13379
rect 27261 13345 27295 13379
rect 6469 13277 6503 13311
rect 7021 13277 7055 13311
rect 10057 13277 10091 13311
rect 14105 13277 14139 13311
rect 14289 13277 14323 13311
rect 15025 13277 15059 13311
rect 15485 13277 15519 13311
rect 15577 13277 15611 13311
rect 15945 13277 15979 13311
rect 16957 13277 16991 13311
rect 17104 13277 17138 13311
rect 18153 13277 18187 13311
rect 19441 13277 19475 13311
rect 19809 13277 19843 13311
rect 23673 13277 23707 13311
rect 23857 13277 23891 13311
rect 24409 13277 24443 13311
rect 25605 13277 25639 13311
rect 25789 13277 25823 13311
rect 26249 13277 26283 13311
rect 26985 13277 27019 13311
rect 27721 13277 27755 13311
rect 27905 13277 27939 13311
rect 30481 13277 30515 13311
rect 31125 13277 31159 13311
rect 31769 13277 31803 13311
rect 32965 13277 32999 13311
rect 33609 13277 33643 13311
rect 34713 13277 34747 13311
rect 7288 13209 7322 13243
rect 8953 13209 8987 13243
rect 9137 13209 9171 13243
rect 10324 13209 10358 13243
rect 12348 13209 12382 13243
rect 16221 13209 16255 13243
rect 24685 13209 24719 13243
rect 27261 13209 27295 13243
rect 34958 13209 34992 13243
rect 11437 13141 11471 13175
rect 25697 13141 25731 13175
rect 30297 13141 30331 13175
rect 31585 13141 31619 13175
rect 36093 13141 36127 13175
rect 4077 12937 4111 12971
rect 9413 12937 9447 12971
rect 20085 12937 20119 12971
rect 2964 12869 2998 12903
rect 7656 12869 7690 12903
rect 9321 12869 9355 12903
rect 12909 12869 12943 12903
rect 17417 12869 17451 12903
rect 18153 12869 18187 12903
rect 19349 12869 19383 12903
rect 19993 12869 20027 12903
rect 30196 12869 30230 12903
rect 32597 12869 32631 12903
rect 2697 12801 2731 12835
rect 7389 12801 7423 12835
rect 10425 12801 10459 12835
rect 12817 12801 12851 12835
rect 13001 12801 13035 12835
rect 14933 12801 14967 12835
rect 15209 12801 15243 12835
rect 16681 12801 16715 12835
rect 16957 12801 16991 12835
rect 18061 12801 18095 12835
rect 18245 12801 18279 12835
rect 18429 12801 18463 12835
rect 18521 12801 18555 12835
rect 19165 12801 19199 12835
rect 19441 12801 19475 12835
rect 20637 12801 20671 12835
rect 20821 12801 20855 12835
rect 23673 12801 23707 12835
rect 23857 12801 23891 12835
rect 28273 12801 28307 12835
rect 28457 12801 28491 12835
rect 28917 12801 28951 12835
rect 29101 12801 29135 12835
rect 32781 12801 32815 12835
rect 10057 12733 10091 12767
rect 10241 12733 10275 12767
rect 11529 12733 11563 12767
rect 11805 12733 11839 12767
rect 18981 12733 19015 12767
rect 29929 12733 29963 12767
rect 8769 12665 8803 12699
rect 10333 12665 10367 12699
rect 15485 12665 15519 12699
rect 16773 12665 16807 12699
rect 17877 12665 17911 12699
rect 10241 12597 10275 12631
rect 15301 12597 15335 12631
rect 20729 12597 20763 12631
rect 23673 12597 23707 12631
rect 28273 12597 28307 12631
rect 28917 12597 28951 12631
rect 31309 12597 31343 12631
rect 32965 12597 32999 12631
rect 8401 12393 8435 12427
rect 10333 12393 10367 12427
rect 14289 12393 14323 12427
rect 14381 12393 14415 12427
rect 16313 12393 16347 12427
rect 17509 12393 17543 12427
rect 19809 12393 19843 12427
rect 22937 12393 22971 12427
rect 26985 12393 27019 12427
rect 30941 12393 30975 12427
rect 15669 12325 15703 12359
rect 17003 12325 17037 12359
rect 17141 12325 17175 12359
rect 18245 12325 18279 12359
rect 29561 12325 29595 12359
rect 7021 12257 7055 12291
rect 14289 12257 14323 12291
rect 17233 12257 17267 12291
rect 22937 12257 22971 12291
rect 23029 12257 23063 12291
rect 27537 12257 27571 12291
rect 9781 12189 9815 12223
rect 10241 12189 10275 12223
rect 10425 12189 10459 12223
rect 14473 12189 14507 12223
rect 15301 12189 15335 12223
rect 16129 12189 16163 12223
rect 18061 12189 18095 12223
rect 20453 12189 20487 12223
rect 23121 12189 23155 12223
rect 23581 12189 23615 12223
rect 23765 12189 23799 12223
rect 24961 12189 24995 12223
rect 25145 12189 25179 12223
rect 25605 12189 25639 12223
rect 25861 12189 25895 12223
rect 27813 12189 27847 12223
rect 28825 12189 28859 12223
rect 29009 12189 29043 12223
rect 29561 12189 29595 12223
rect 29745 12189 29779 12223
rect 30757 12189 30791 12223
rect 31769 12189 31803 12223
rect 33425 12189 33459 12223
rect 7288 12121 7322 12155
rect 14105 12121 14139 12155
rect 15485 12121 15519 12155
rect 16865 12121 16899 12155
rect 19717 12121 19751 12155
rect 20720 12121 20754 12155
rect 22753 12121 22787 12155
rect 30573 12121 30607 12155
rect 32597 12121 32631 12155
rect 32781 12121 32815 12155
rect 33609 12121 33643 12155
rect 9597 12053 9631 12087
rect 21833 12053 21867 12087
rect 23765 12053 23799 12087
rect 25053 12053 25087 12087
rect 28917 12053 28951 12087
rect 31585 12053 31619 12087
rect 32965 12053 32999 12087
rect 33793 12053 33827 12087
rect 7941 11849 7975 11883
rect 13553 11849 13587 11883
rect 17325 11849 17359 11883
rect 19073 11849 19107 11883
rect 23213 11849 23247 11883
rect 25145 11849 25179 11883
rect 34069 11849 34103 11883
rect 14381 11781 14415 11815
rect 16865 11781 16899 11815
rect 19695 11781 19729 11815
rect 24032 11781 24066 11815
rect 8125 11713 8159 11747
rect 12633 11713 12667 11747
rect 13461 11713 13495 11747
rect 17141 11713 17175 11747
rect 18889 11713 18923 11747
rect 19993 11713 20027 11747
rect 21097 11713 21131 11747
rect 21281 11713 21315 11747
rect 21833 11713 21867 11747
rect 22089 11713 22123 11747
rect 23765 11713 23799 11747
rect 25605 11713 25639 11747
rect 25789 11713 25823 11747
rect 26985 11713 27019 11747
rect 27169 11713 27203 11747
rect 28365 11713 28399 11747
rect 28549 11713 28583 11747
rect 31585 11713 31619 11747
rect 32945 11713 32979 11747
rect 34713 11713 34747 11747
rect 12909 11645 12943 11679
rect 16129 11645 16163 11679
rect 16957 11645 16991 11679
rect 19809 11645 19843 11679
rect 21189 11645 21223 11679
rect 28733 11645 28767 11679
rect 32689 11645 32723 11679
rect 19625 11577 19659 11611
rect 19901 11577 19935 11611
rect 31401 11577 31435 11611
rect 12449 11509 12483 11543
rect 12817 11509 12851 11543
rect 16865 11509 16899 11543
rect 25697 11509 25731 11543
rect 26985 11509 27019 11543
rect 34529 11509 34563 11543
rect 15577 11305 15611 11339
rect 18061 11305 18095 11339
rect 18429 11305 18463 11339
rect 20637 11305 20671 11339
rect 21373 11305 21407 11339
rect 21465 11305 21499 11339
rect 25789 11305 25823 11339
rect 28549 11305 28583 11339
rect 13461 11237 13495 11271
rect 16405 11237 16439 11271
rect 17233 11237 17267 11271
rect 17417 11237 17451 11271
rect 33701 11237 33735 11271
rect 14749 11169 14783 11203
rect 16957 11169 16991 11203
rect 23305 11169 23339 11203
rect 30021 11169 30055 11203
rect 9965 11101 9999 11135
rect 10149 11101 10183 11135
rect 12081 11101 12115 11135
rect 12348 11101 12382 11135
rect 14565 11101 14599 11135
rect 17969 11101 18003 11135
rect 19257 11101 19291 11135
rect 21189 11101 21223 11135
rect 21327 11101 21361 11135
rect 21557 11101 21591 11135
rect 23029 11101 23063 11135
rect 24409 11101 24443 11135
rect 27169 11101 27203 11135
rect 32413 11101 32447 11135
rect 14381 11033 14415 11067
rect 15209 11033 15243 11067
rect 15393 11033 15427 11067
rect 16037 11033 16071 11067
rect 16221 11033 16255 11067
rect 19524 11033 19558 11067
rect 24676 11033 24710 11067
rect 27436 11033 27470 11067
rect 30288 11033 30322 11067
rect 10057 10965 10091 10999
rect 31401 10965 31435 10999
rect 14565 10761 14599 10795
rect 17141 10761 17175 10795
rect 20085 10761 20119 10795
rect 34069 10761 34103 10795
rect 16129 10693 16163 10727
rect 19165 10693 19199 10727
rect 24225 10693 24259 10727
rect 24777 10693 24811 10727
rect 30735 10693 30769 10727
rect 32956 10693 32990 10727
rect 8677 10625 8711 10659
rect 8944 10625 8978 10659
rect 10977 10625 11011 10659
rect 11529 10625 11563 10659
rect 11785 10625 11819 10659
rect 14013 10625 14047 10659
rect 15117 10625 15151 10659
rect 15577 10625 15611 10659
rect 15945 10625 15979 10659
rect 16681 10625 16715 10659
rect 16773 10625 16807 10659
rect 16957 10625 16991 10659
rect 19533 10625 19567 10659
rect 19993 10625 20027 10659
rect 20177 10625 20211 10659
rect 24041 10625 24075 10659
rect 25145 10625 25179 10659
rect 27675 10625 27709 10659
rect 27905 10625 27939 10659
rect 29423 10625 29457 10659
rect 29653 10625 29687 10659
rect 31033 10625 31067 10659
rect 10793 10557 10827 10591
rect 14289 10557 14323 10591
rect 19349 10557 19383 10591
rect 24961 10557 24995 10591
rect 27813 10557 27847 10591
rect 30849 10557 30883 10591
rect 32689 10557 32723 10591
rect 10057 10489 10091 10523
rect 10609 10489 10643 10523
rect 10885 10489 10919 10523
rect 12909 10489 12943 10523
rect 27537 10489 27571 10523
rect 29285 10489 29319 10523
rect 30665 10489 30699 10523
rect 10793 10421 10827 10455
rect 14105 10421 14139 10455
rect 19349 10421 19383 10455
rect 19441 10421 19475 10455
rect 24961 10421 24995 10455
rect 25053 10421 25087 10455
rect 27721 10421 27755 10455
rect 29469 10421 29503 10455
rect 29561 10421 29595 10455
rect 30941 10421 30975 10455
rect 10977 10217 11011 10251
rect 14657 10217 14691 10251
rect 15025 10217 15059 10251
rect 16497 10217 16531 10251
rect 18613 10217 18647 10251
rect 26985 10217 27019 10251
rect 27537 10217 27571 10251
rect 30941 10217 30975 10251
rect 34069 10217 34103 10251
rect 15761 10149 15795 10183
rect 10793 10081 10827 10115
rect 14749 10081 14783 10115
rect 29561 10081 29595 10115
rect 29837 10081 29871 10115
rect 1869 10013 1903 10047
rect 9137 10013 9171 10047
rect 11253 10013 11287 10047
rect 12633 10013 12667 10047
rect 12817 10013 12851 10047
rect 14657 10013 14691 10047
rect 15577 10013 15611 10047
rect 17233 10013 17267 10047
rect 20545 10013 20579 10047
rect 24869 10013 24903 10047
rect 25605 10013 25639 10047
rect 27445 10013 27479 10047
rect 27629 10013 27663 10047
rect 28825 10013 28859 10047
rect 29009 10013 29043 10047
rect 30849 10013 30883 10047
rect 31033 10013 31067 10047
rect 32229 10013 32263 10047
rect 32689 10013 32723 10047
rect 12909 9945 12943 9979
rect 16221 9945 16255 9979
rect 16405 9945 16439 9979
rect 17500 9945 17534 9979
rect 20812 9945 20846 9979
rect 25872 9945 25906 9979
rect 32934 9945 32968 9979
rect 1961 9877 1995 9911
rect 8953 9877 8987 9911
rect 11161 9877 11195 9911
rect 21925 9877 21959 9911
rect 24961 9877 24995 9911
rect 28917 9877 28951 9911
rect 32045 9877 32079 9911
rect 17509 9673 17543 9707
rect 20913 9673 20947 9707
rect 25329 9673 25363 9707
rect 26157 9673 26191 9707
rect 29929 9673 29963 9707
rect 8208 9605 8242 9639
rect 15209 9605 15243 9639
rect 19809 9605 19843 9639
rect 25237 9605 25271 9639
rect 28816 9605 28850 9639
rect 30849 9605 30883 9639
rect 10333 9537 10367 9571
rect 11989 9537 12023 9571
rect 13093 9537 13127 9571
rect 15025 9537 15059 9571
rect 17693 9537 17727 9571
rect 19165 9537 19199 9571
rect 21097 9537 21131 9571
rect 21925 9537 21959 9571
rect 22192 9537 22226 9571
rect 24501 9537 24535 9571
rect 26065 9537 26099 9571
rect 26249 9537 26283 9571
rect 26985 9537 27019 9571
rect 27353 9537 27387 9571
rect 31217 9537 31251 9571
rect 32137 9537 32171 9571
rect 32321 9537 32355 9571
rect 7941 9469 7975 9503
rect 13369 9469 13403 9503
rect 24317 9469 24351 9503
rect 27169 9469 27203 9503
rect 28549 9469 28583 9503
rect 31033 9469 31067 9503
rect 31125 9469 31159 9503
rect 9321 9401 9355 9435
rect 19993 9401 20027 9435
rect 10149 9333 10183 9367
rect 11805 9333 11839 9367
rect 12909 9333 12943 9367
rect 13277 9333 13311 9367
rect 18981 9333 19015 9367
rect 23305 9333 23339 9367
rect 24685 9333 24719 9367
rect 27169 9333 27203 9367
rect 27261 9333 27295 9367
rect 31033 9333 31067 9367
rect 32229 9333 32263 9367
rect 9321 9129 9355 9163
rect 16221 9129 16255 9163
rect 18705 9129 18739 9163
rect 21557 9129 21591 9163
rect 33149 9129 33183 9163
rect 13093 9061 13127 9095
rect 16589 9061 16623 9095
rect 11713 8993 11747 9027
rect 17325 8993 17359 9027
rect 18337 8993 18371 9027
rect 27629 8993 27663 9027
rect 8953 8925 8987 8959
rect 9137 8925 9171 8959
rect 9781 8925 9815 8959
rect 11969 8925 12003 8959
rect 14657 8925 14691 8959
rect 14841 8925 14875 8959
rect 15025 8925 15059 8959
rect 15669 8925 15703 8959
rect 16129 8925 16163 8959
rect 17049 8925 17083 8959
rect 18521 8925 18555 8959
rect 19257 8925 19291 8959
rect 19513 8925 19547 8959
rect 21189 8925 21223 8959
rect 21373 8925 21407 8959
rect 22063 8925 22097 8959
rect 22385 8925 22419 8959
rect 23029 8925 23063 8959
rect 23305 8925 23339 8959
rect 24409 8925 24443 8959
rect 27813 8925 27847 8959
rect 31033 8925 31067 8959
rect 10048 8857 10082 8891
rect 22201 8857 22235 8891
rect 22293 8857 22327 8891
rect 24676 8857 24710 8891
rect 31300 8857 31334 8891
rect 33057 8857 33091 8891
rect 11161 8789 11195 8823
rect 15485 8789 15519 8823
rect 20637 8789 20671 8823
rect 22569 8789 22603 8823
rect 25789 8789 25823 8823
rect 27997 8789 28031 8823
rect 32413 8789 32447 8823
rect 8769 8585 8803 8619
rect 14105 8585 14139 8619
rect 18061 8585 18095 8619
rect 19533 8585 19567 8619
rect 24961 8585 24995 8619
rect 25605 8585 25639 8619
rect 8493 8517 8527 8551
rect 10977 8517 11011 8551
rect 18797 8517 18831 8551
rect 22201 8517 22235 8551
rect 24593 8517 24627 8551
rect 24685 8517 24719 8551
rect 7665 8449 7699 8483
rect 8217 8449 8251 8483
rect 8401 8449 8435 8483
rect 8585 8449 8619 8483
rect 9229 8449 9263 8483
rect 11529 8449 11563 8483
rect 11713 8449 11747 8483
rect 11805 8449 11839 8483
rect 11943 8449 11977 8483
rect 12725 8449 12759 8483
rect 12992 8449 13026 8483
rect 14657 8449 14691 8483
rect 14924 8449 14958 8483
rect 17509 8449 17543 8483
rect 17693 8449 17727 8483
rect 17785 8449 17819 8483
rect 17923 8449 17957 8483
rect 18521 8449 18555 8483
rect 18705 8449 18739 8483
rect 18935 8449 18969 8483
rect 19717 8449 19751 8483
rect 24409 8449 24443 8483
rect 24777 8449 24811 8483
rect 25421 8449 25455 8483
rect 26433 8449 26467 8483
rect 26985 8449 27019 8483
rect 27241 8449 27275 8483
rect 29469 8449 29503 8483
rect 29653 8449 29687 8483
rect 32853 8449 32887 8483
rect 34621 8449 34655 8483
rect 34805 8449 34839 8483
rect 20177 8381 20211 8415
rect 20453 8381 20487 8415
rect 32597 8381 32631 8415
rect 16037 8313 16071 8347
rect 23489 8313 23523 8347
rect 26249 8313 26283 8347
rect 28365 8313 28399 8347
rect 33977 8313 34011 8347
rect 7481 8245 7515 8279
rect 12081 8245 12115 8279
rect 19073 8245 19107 8279
rect 29837 8245 29871 8279
rect 34989 8245 35023 8279
rect 8217 8041 8251 8075
rect 11069 8041 11103 8075
rect 11989 8041 12023 8075
rect 15025 8041 15059 8075
rect 18705 8041 18739 8075
rect 21189 8041 21223 8075
rect 21649 8041 21683 8075
rect 25145 8041 25179 8075
rect 28917 8041 28951 8075
rect 31309 8041 31343 8075
rect 33057 8041 33091 8075
rect 33149 8041 33183 8075
rect 15577 7973 15611 8007
rect 16681 7973 16715 8007
rect 23397 7973 23431 8007
rect 32321 7973 32355 8007
rect 10701 7905 10735 7939
rect 11621 7905 11655 7939
rect 16313 7905 16347 7939
rect 16773 7905 16807 7939
rect 18337 7905 18371 7939
rect 19901 7905 19935 7939
rect 22661 7905 22695 7939
rect 32873 7905 32907 7939
rect 33057 7905 33091 7939
rect 34713 7905 34747 7939
rect 6837 7837 6871 7871
rect 9689 7837 9723 7871
rect 9873 7837 9907 7871
rect 10057 7837 10091 7871
rect 10885 7837 10919 7871
rect 11805 7837 11839 7871
rect 14473 7837 14507 7871
rect 14657 7837 14691 7871
rect 14841 7837 14875 7871
rect 15485 7837 15519 7871
rect 18521 7837 18555 7871
rect 20637 7837 20671 7871
rect 21005 7837 21039 7871
rect 21833 7837 21867 7871
rect 22293 7837 22327 7871
rect 22477 7837 22511 7871
rect 23213 7837 23247 7871
rect 24409 7837 24443 7871
rect 25329 7837 25363 7871
rect 26525 7837 26559 7871
rect 26893 7837 26927 7871
rect 27537 7837 27571 7871
rect 29929 7837 29963 7871
rect 32229 7837 32263 7871
rect 32413 7837 32447 7871
rect 33241 7837 33275 7871
rect 34161 7837 34195 7871
rect 7104 7769 7138 7803
rect 9965 7769 9999 7803
rect 14749 7769 14783 7803
rect 17693 7769 17727 7803
rect 19717 7769 19751 7803
rect 20821 7769 20855 7803
rect 20913 7769 20947 7803
rect 26709 7769 26743 7803
rect 26801 7769 26835 7803
rect 27804 7769 27838 7803
rect 30174 7769 30208 7803
rect 34958 7769 34992 7803
rect 10241 7701 10275 7735
rect 17785 7701 17819 7735
rect 24593 7701 24627 7735
rect 27077 7701 27111 7735
rect 33977 7701 34011 7735
rect 36093 7701 36127 7735
rect 9413 7497 9447 7531
rect 14933 7497 14967 7531
rect 18337 7497 18371 7531
rect 35173 7497 35207 7531
rect 8217 7429 8251 7463
rect 13001 7429 13035 7463
rect 13093 7429 13127 7463
rect 15669 7429 15703 7463
rect 19717 7429 19751 7463
rect 21281 7429 21315 7463
rect 23121 7429 23155 7463
rect 23305 7429 23339 7463
rect 23857 7429 23891 7463
rect 27353 7429 27387 7463
rect 28641 7429 28675 7463
rect 28733 7429 28767 7463
rect 34897 7429 34931 7463
rect 8033 7361 8067 7395
rect 8309 7361 8343 7395
rect 8401 7361 8435 7395
rect 9229 7361 9263 7395
rect 12725 7361 12759 7395
rect 13809 7361 13843 7395
rect 15485 7361 15519 7395
rect 17141 7361 17175 7395
rect 18153 7361 18187 7395
rect 18981 7361 19015 7395
rect 20545 7361 20579 7395
rect 21097 7361 21131 7395
rect 22385 7361 22419 7395
rect 23765 7361 23799 7395
rect 23949 7361 23983 7395
rect 26341 7361 26375 7395
rect 27169 7361 27203 7395
rect 27997 7361 28031 7395
rect 28457 7361 28491 7395
rect 28825 7361 28859 7395
rect 29653 7361 29687 7395
rect 30380 7361 30414 7395
rect 32597 7361 32631 7395
rect 32781 7361 32815 7395
rect 34621 7361 34655 7395
rect 34805 7361 34839 7395
rect 34989 7361 35023 7395
rect 9045 7293 9079 7327
rect 12633 7293 12667 7327
rect 13553 7293 13587 7327
rect 19901 7293 19935 7327
rect 22201 7293 22235 7327
rect 24869 7293 24903 7327
rect 25145 7293 25179 7327
rect 26985 7293 27019 7327
rect 30113 7293 30147 7327
rect 8585 7225 8619 7259
rect 19165 7225 19199 7259
rect 12449 7157 12483 7191
rect 17233 7157 17267 7191
rect 20361 7157 20395 7191
rect 22569 7157 22603 7191
rect 26157 7157 26191 7191
rect 27813 7157 27847 7191
rect 29009 7157 29043 7191
rect 29469 7157 29503 7191
rect 31493 7157 31527 7191
rect 32689 7157 32723 7191
rect 18061 6953 18095 6987
rect 19717 6953 19751 6987
rect 27721 6953 27755 6987
rect 34713 6953 34747 6987
rect 21649 6885 21683 6919
rect 9873 6817 9907 6851
rect 13461 6817 13495 6851
rect 16129 6817 16163 6851
rect 22385 6817 22419 6851
rect 34897 6817 34931 6851
rect 9229 6749 9263 6783
rect 9413 6749 9447 6783
rect 11713 6749 11747 6783
rect 11897 6749 11931 6783
rect 12081 6749 12115 6783
rect 12725 6749 12759 6783
rect 13369 6749 13403 6783
rect 13553 6749 13587 6783
rect 15485 6749 15519 6783
rect 15669 6749 15703 6783
rect 18061 6749 18095 6783
rect 18245 6749 18279 6783
rect 19533 6749 19567 6783
rect 20269 6749 20303 6783
rect 24593 6749 24627 6783
rect 25237 6749 25271 6783
rect 25881 6749 25915 6783
rect 26433 6749 26467 6783
rect 28825 6749 28859 6783
rect 29561 6749 29595 6783
rect 29929 6749 29963 6783
rect 30573 6749 30607 6783
rect 30757 6749 30791 6783
rect 31769 6749 31803 6783
rect 32413 6749 32447 6783
rect 32680 6749 32714 6783
rect 34989 6749 35023 6783
rect 10118 6681 10152 6715
rect 15577 6681 15611 6715
rect 16374 6681 16408 6715
rect 20514 6681 20548 6715
rect 22652 6681 22686 6715
rect 29745 6681 29779 6715
rect 29837 6681 29871 6715
rect 34713 6681 34747 6715
rect 11253 6613 11287 6647
rect 12541 6613 12575 6647
rect 17509 6613 17543 6647
rect 23765 6613 23799 6647
rect 24409 6613 24443 6647
rect 25053 6613 25087 6647
rect 25697 6613 25731 6647
rect 28641 6613 28675 6647
rect 30113 6613 30147 6647
rect 30941 6613 30975 6647
rect 31585 6613 31619 6647
rect 33793 6613 33827 6647
rect 35173 6613 35207 6647
rect 9781 6409 9815 6443
rect 13553 6409 13587 6443
rect 14197 6409 14231 6443
rect 15117 6409 15151 6443
rect 17509 6409 17543 6443
rect 20361 6409 20395 6443
rect 22385 6409 22419 6443
rect 22845 6409 22879 6443
rect 24501 6409 24535 6443
rect 26433 6409 26467 6443
rect 28089 6409 28123 6443
rect 29745 6409 29779 6443
rect 30297 6409 30331 6443
rect 30941 6409 30975 6443
rect 33885 6409 33919 6443
rect 10701 6341 10735 6375
rect 11980 6341 12014 6375
rect 16751 6341 16785 6375
rect 18797 6341 18831 6375
rect 24409 6341 24443 6375
rect 32229 6341 32263 6375
rect 33057 6341 33091 6375
rect 7757 6273 7791 6307
rect 7941 6273 7975 6307
rect 8401 6273 8435 6307
rect 8657 6273 8691 6307
rect 10425 6273 10459 6307
rect 10609 6273 10643 6307
rect 10793 6273 10827 6307
rect 13737 6273 13771 6307
rect 14381 6273 14415 6307
rect 15301 6273 15335 6307
rect 17049 6273 17083 6307
rect 17693 6273 17727 6307
rect 18521 6273 18555 6307
rect 18705 6273 18739 6307
rect 18889 6273 18923 6307
rect 20085 6273 20119 6307
rect 20177 6273 20211 6307
rect 21097 6273 21131 6307
rect 21833 6273 21867 6307
rect 22017 6273 22051 6307
rect 22109 6273 22143 6307
rect 22201 6273 22235 6307
rect 23029 6273 23063 6307
rect 23765 6273 23799 6307
rect 25053 6273 25087 6307
rect 25320 6273 25354 6307
rect 27077 6273 27111 6307
rect 27261 6273 27295 6307
rect 27353 6273 27387 6307
rect 27445 6273 27479 6307
rect 28273 6273 28307 6307
rect 29193 6273 29227 6307
rect 29331 6273 29365 6307
rect 29469 6273 29503 6307
rect 29561 6273 29595 6307
rect 30481 6273 30515 6307
rect 31125 6273 31159 6307
rect 32597 6273 32631 6307
rect 33425 6273 33459 6307
rect 34069 6273 34103 6307
rect 7849 6205 7883 6239
rect 11713 6205 11747 6239
rect 16681 6205 16715 6239
rect 16865 6205 16899 6239
rect 32299 6205 32333 6239
rect 32413 6205 32447 6239
rect 33241 6205 33275 6239
rect 16957 6137 16991 6171
rect 19073 6137 19107 6171
rect 32505 6137 32539 6171
rect 33333 6137 33367 6171
rect 10977 6069 11011 6103
rect 13093 6069 13127 6103
rect 21189 6069 21223 6103
rect 23581 6069 23615 6103
rect 27629 6069 27663 6103
rect 33241 6069 33275 6103
rect 9137 5865 9171 5899
rect 9965 5865 9999 5899
rect 17785 5865 17819 5899
rect 21741 5865 21775 5899
rect 26709 5865 26743 5899
rect 28549 5865 28583 5899
rect 28641 5865 28675 5899
rect 30849 5865 30883 5899
rect 36093 5865 36127 5899
rect 37933 5865 37967 5899
rect 9229 5797 9263 5831
rect 17141 5797 17175 5831
rect 29561 5797 29595 5831
rect 30205 5797 30239 5831
rect 31493 5797 31527 5831
rect 9137 5729 9171 5763
rect 10977 5729 11011 5763
rect 13001 5729 13035 5763
rect 19257 5729 19291 5763
rect 25329 5729 25363 5763
rect 28549 5729 28583 5763
rect 9321 5661 9355 5695
rect 10149 5661 10183 5695
rect 10609 5661 10643 5695
rect 10793 5661 10827 5695
rect 11437 5661 11471 5695
rect 11621 5661 11655 5695
rect 11805 5661 11839 5695
rect 12725 5661 12759 5695
rect 14657 5661 14691 5695
rect 16681 5661 16715 5695
rect 17325 5661 17359 5695
rect 17969 5661 18003 5695
rect 18705 5661 18739 5695
rect 22385 5661 22419 5695
rect 23673 5661 23707 5695
rect 24409 5661 24443 5695
rect 24593 5661 24627 5695
rect 25053 5661 25087 5695
rect 26341 5661 26375 5695
rect 26525 5661 26559 5695
rect 27353 5661 27387 5695
rect 28733 5661 28767 5695
rect 29745 5661 29779 5695
rect 30389 5661 30423 5695
rect 31033 5661 31067 5695
rect 31677 5661 31711 5695
rect 32321 5661 32355 5695
rect 34713 5661 34747 5695
rect 38117 5661 38151 5695
rect 8953 5593 8987 5627
rect 11713 5593 11747 5627
rect 14924 5593 14958 5627
rect 19502 5593 19536 5627
rect 21649 5593 21683 5627
rect 23857 5593 23891 5627
rect 28365 5593 28399 5627
rect 34958 5593 34992 5627
rect 11989 5525 12023 5559
rect 16037 5525 16071 5559
rect 16497 5525 16531 5559
rect 18521 5525 18555 5559
rect 20637 5525 20671 5559
rect 22477 5525 22511 5559
rect 24501 5525 24535 5559
rect 27169 5525 27203 5559
rect 33609 5525 33643 5559
rect 9505 5321 9539 5355
rect 10609 5321 10643 5355
rect 11713 5321 11747 5355
rect 18705 5321 18739 5355
rect 26433 5321 26467 5355
rect 31585 5321 31619 5355
rect 34437 5321 34471 5355
rect 14381 5253 14415 5287
rect 21005 5253 21039 5287
rect 27230 5253 27264 5287
rect 32382 5253 32416 5287
rect 9689 5185 9723 5219
rect 10793 5185 10827 5219
rect 11897 5185 11931 5219
rect 12808 5185 12842 5219
rect 17233 5185 17267 5219
rect 17417 5185 17451 5219
rect 18245 5185 18279 5219
rect 18889 5185 18923 5219
rect 19419 5185 19453 5219
rect 19717 5185 19751 5219
rect 20453 5185 20487 5219
rect 22017 5185 22051 5219
rect 22753 5185 22787 5219
rect 23397 5185 23431 5219
rect 23664 5185 23698 5219
rect 25329 5185 25363 5219
rect 26249 5185 26283 5219
rect 26433 5185 26467 5219
rect 28825 5185 28859 5219
rect 29081 5185 29115 5219
rect 30665 5185 30699 5219
rect 30849 5185 30883 5219
rect 31401 5185 31435 5219
rect 31585 5185 31619 5219
rect 34621 5185 34655 5219
rect 35265 5185 35299 5219
rect 37841 5185 37875 5219
rect 12541 5117 12575 5151
rect 16129 5117 16163 5151
rect 19533 5117 19567 5151
rect 26985 5117 27019 5151
rect 32137 5117 32171 5151
rect 19349 5049 19383 5083
rect 20269 5049 20303 5083
rect 21833 5049 21867 5083
rect 35081 5049 35115 5083
rect 13921 4981 13955 5015
rect 17325 4981 17359 5015
rect 18061 4981 18095 5015
rect 19625 4981 19659 5015
rect 21097 4981 21131 5015
rect 22845 4981 22879 5015
rect 24777 4981 24811 5015
rect 25421 4981 25455 5015
rect 28365 4981 28399 5015
rect 30205 4981 30239 5015
rect 30757 4981 30791 5015
rect 33517 4981 33551 5015
rect 38025 4981 38059 5015
rect 14289 4777 14323 4811
rect 14381 4777 14415 4811
rect 15577 4777 15611 4811
rect 19349 4777 19383 4811
rect 22017 4777 22051 4811
rect 24593 4777 24627 4811
rect 24685 4777 24719 4811
rect 26617 4777 26651 4811
rect 26709 4777 26743 4811
rect 27997 4777 28031 4811
rect 28825 4777 28859 4811
rect 32413 4777 32447 4811
rect 33609 4777 33643 4811
rect 35725 4777 35759 4811
rect 37197 4777 37231 4811
rect 10241 4709 10275 4743
rect 14105 4709 14139 4743
rect 15371 4709 15405 4743
rect 27261 4709 27295 4743
rect 32873 4709 32907 4743
rect 14289 4641 14323 4675
rect 15485 4641 15519 4675
rect 16221 4641 16255 4675
rect 21741 4641 21775 4675
rect 21879 4641 21913 4675
rect 24409 4641 24443 4675
rect 24593 4641 24627 4675
rect 26433 4641 26467 4675
rect 26617 4641 26651 4675
rect 32505 4641 32539 4675
rect 9045 4573 9079 4607
rect 9229 4573 9263 4607
rect 10425 4573 10459 4607
rect 11529 4573 11563 4607
rect 12265 4573 12299 4607
rect 12909 4573 12943 4607
rect 13553 4573 13587 4607
rect 14473 4573 14507 4607
rect 15669 4573 15703 4607
rect 16129 4573 16163 4607
rect 16313 4573 16347 4607
rect 16865 4573 16899 4607
rect 19257 4573 19291 4607
rect 19441 4573 19475 4607
rect 20085 4573 20119 4607
rect 21097 4573 21131 4607
rect 21281 4573 21315 4607
rect 22109 4573 22143 4607
rect 22569 4573 22603 4607
rect 23305 4573 23339 4607
rect 24777 4573 24811 4607
rect 25605 4573 25639 4607
rect 26801 4573 26835 4607
rect 27445 4573 27479 4607
rect 27905 4573 27939 4607
rect 28089 4573 28123 4607
rect 28733 4573 28767 4607
rect 28825 4573 28859 4607
rect 30113 4573 30147 4607
rect 32689 4573 32723 4607
rect 33793 4573 33827 4607
rect 34713 4573 34747 4607
rect 35081 4573 35115 4607
rect 35909 4573 35943 4607
rect 37381 4573 37415 4607
rect 37841 4573 37875 4607
rect 15301 4505 15335 4539
rect 17132 4505 17166 4539
rect 21811 4505 21845 4539
rect 28549 4505 28583 4539
rect 30380 4505 30414 4539
rect 32413 4505 32447 4539
rect 34897 4505 34931 4539
rect 34989 4505 35023 4539
rect 9137 4437 9171 4471
rect 11345 4437 11379 4471
rect 12081 4437 12115 4471
rect 12725 4437 12759 4471
rect 13369 4437 13403 4471
rect 18245 4437 18279 4471
rect 19901 4437 19935 4471
rect 21281 4437 21315 4471
rect 22753 4437 22787 4471
rect 23489 4437 23523 4471
rect 25421 4437 25455 4471
rect 29009 4437 29043 4471
rect 31493 4437 31527 4471
rect 35265 4437 35299 4471
rect 38025 4437 38059 4471
rect 11989 4233 12023 4267
rect 19441 4233 19475 4267
rect 23213 4233 23247 4267
rect 34713 4233 34747 4267
rect 36553 4233 36587 4267
rect 8852 4165 8886 4199
rect 11529 4165 11563 4199
rect 12817 4165 12851 4199
rect 15393 4165 15427 4199
rect 18981 4165 19015 4199
rect 20269 4165 20303 4199
rect 22100 4165 22134 4199
rect 24041 4165 24075 4199
rect 29377 4165 29411 4199
rect 30573 4165 30607 4199
rect 8585 4097 8619 4131
rect 10793 4097 10827 4131
rect 11805 4097 11839 4131
rect 12541 4097 12575 4131
rect 12725 4097 12759 4131
rect 12909 4097 12943 4131
rect 13921 4097 13955 4131
rect 14105 4097 14139 4131
rect 14657 4097 14691 4131
rect 15669 4097 15703 4131
rect 16865 4097 16899 4131
rect 17325 4097 17359 4131
rect 17693 4097 17727 4131
rect 18337 4097 18371 4131
rect 19257 4097 19291 4131
rect 21097 4097 21131 4131
rect 24961 4097 24995 4131
rect 25973 4097 26007 4131
rect 26985 4097 27019 4131
rect 27721 4097 27755 4131
rect 28641 4097 28675 4131
rect 29653 4097 29687 4131
rect 30941 4097 30975 4131
rect 31585 4097 31619 4131
rect 32321 4097 32355 4131
rect 32965 4097 32999 4131
rect 33609 4097 33643 4131
rect 34529 4097 34563 4131
rect 35357 4097 35391 4131
rect 36001 4097 36035 4131
rect 36737 4097 36771 4131
rect 37657 4097 37691 4131
rect 10609 4029 10643 4063
rect 10701 4029 10735 4063
rect 11621 4029 11655 4063
rect 14013 4029 14047 4063
rect 15485 4029 15519 4063
rect 17509 4029 17543 4063
rect 19165 4029 19199 4063
rect 21833 4029 21867 4063
rect 24685 4029 24719 4063
rect 29469 4029 29503 4063
rect 30757 4029 30791 4063
rect 30849 4029 30883 4063
rect 34345 4029 34379 4063
rect 9965 3961 9999 3995
rect 10425 3961 10459 3995
rect 15853 3961 15887 3995
rect 17601 3961 17635 3995
rect 24225 3961 24259 3995
rect 28457 3961 28491 3995
rect 32781 3961 32815 3995
rect 35817 3961 35851 3995
rect 1961 3893 1995 3927
rect 10609 3893 10643 3927
rect 11529 3893 11563 3927
rect 13093 3893 13127 3927
rect 14841 3893 14875 3927
rect 15485 3893 15519 3927
rect 16681 3893 16715 3927
rect 17509 3893 17543 3927
rect 18153 3893 18187 3927
rect 19257 3893 19291 3927
rect 20361 3893 20395 3927
rect 20913 3893 20947 3927
rect 26157 3893 26191 3927
rect 27169 3893 27203 3927
rect 27905 3893 27939 3927
rect 29653 3893 29687 3927
rect 29837 3893 29871 3927
rect 30757 3893 30791 3927
rect 31401 3893 31435 3927
rect 32137 3893 32171 3927
rect 33425 3893 33459 3927
rect 35173 3893 35207 3927
rect 37841 3893 37875 3927
rect 3801 3689 3835 3723
rect 6561 3689 6595 3723
rect 9137 3689 9171 3723
rect 9229 3689 9263 3723
rect 11161 3689 11195 3723
rect 13001 3689 13035 3723
rect 14473 3689 14507 3723
rect 16865 3689 16899 3723
rect 17325 3689 17359 3723
rect 21373 3689 21407 3723
rect 24593 3689 24627 3723
rect 24961 3689 24995 3723
rect 27169 3689 27203 3723
rect 7573 3621 7607 3655
rect 23857 3621 23891 3655
rect 32873 3621 32907 3655
rect 35265 3621 35299 3655
rect 8953 3553 8987 3587
rect 9137 3553 9171 3587
rect 9770 3553 9804 3587
rect 14105 3553 14139 3587
rect 22477 3553 22511 3587
rect 24593 3553 24627 3587
rect 25881 3553 25915 3587
rect 26157 3553 26191 3587
rect 27813 3553 27847 3587
rect 1593 3485 1627 3519
rect 2697 3485 2731 3519
rect 3985 3485 4019 3519
rect 6745 3485 6779 3519
rect 7757 3485 7791 3519
rect 8217 3485 8251 3519
rect 8401 3485 8435 3519
rect 9321 3485 9355 3519
rect 10048 3485 10082 3519
rect 11621 3485 11655 3519
rect 14289 3485 14323 3519
rect 15485 3485 15519 3519
rect 17509 3485 17543 3519
rect 18521 3485 18555 3519
rect 19993 3485 20027 3519
rect 22017 3485 22051 3519
rect 24501 3485 24535 3519
rect 24777 3485 24811 3519
rect 27353 3485 27387 3519
rect 27997 3485 28031 3519
rect 28181 3485 28215 3519
rect 28825 3485 28859 3519
rect 30021 3485 30055 3519
rect 30113 3485 30147 3519
rect 30757 3485 30791 3519
rect 31861 3485 31895 3519
rect 32045 3485 32079 3519
rect 32137 3485 32171 3519
rect 32229 3485 32263 3519
rect 33057 3485 33091 3519
rect 33793 3485 33827 3519
rect 33977 3485 34011 3519
rect 34713 3485 34747 3519
rect 34989 3485 35023 3519
rect 35081 3485 35115 3519
rect 35725 3485 35759 3519
rect 36553 3485 36587 3519
rect 11888 3417 11922 3451
rect 15752 3417 15786 3451
rect 19349 3417 19383 3451
rect 20260 3417 20294 3451
rect 22722 3417 22756 3451
rect 34897 3417 34931 3451
rect 37933 3417 37967 3451
rect 1409 3349 1443 3383
rect 2513 3349 2547 3383
rect 8309 3349 8343 3383
rect 18337 3349 18371 3383
rect 19441 3349 19475 3383
rect 21833 3349 21867 3383
rect 28641 3349 28675 3383
rect 30297 3349 30331 3383
rect 30941 3349 30975 3383
rect 32413 3349 32447 3383
rect 34161 3349 34195 3383
rect 35909 3349 35943 3383
rect 36737 3349 36771 3383
rect 38025 3349 38059 3383
rect 3065 3145 3099 3179
rect 3801 3145 3835 3179
rect 4629 3145 4663 3179
rect 5181 3145 5215 3179
rect 6377 3145 6411 3179
rect 8953 3145 8987 3179
rect 9965 3145 9999 3179
rect 12909 3145 12943 3179
rect 15485 3145 15519 3179
rect 19257 3145 19291 3179
rect 22937 3145 22971 3179
rect 26433 3145 26467 3179
rect 28733 3145 28767 3179
rect 36553 3145 36587 3179
rect 2881 3077 2915 3111
rect 10977 3077 11011 3111
rect 11713 3077 11747 3111
rect 11805 3077 11839 3111
rect 13706 3077 13740 3111
rect 16957 3077 16991 3111
rect 18144 3077 18178 3111
rect 19993 3077 20027 3111
rect 20913 3077 20947 3111
rect 23857 3077 23891 3111
rect 27620 3077 27654 3111
rect 34244 3077 34278 3111
rect 1409 3009 1443 3043
rect 3985 3009 4019 3043
rect 4813 3009 4847 3043
rect 5457 3009 5491 3043
rect 6561 3009 6595 3043
rect 7573 3009 7607 3043
rect 7840 3009 7874 3043
rect 10149 3009 10183 3043
rect 10793 3009 10827 3043
rect 11529 3009 11563 3043
rect 11897 3009 11931 3043
rect 12541 3009 12575 3043
rect 12725 3009 12759 3043
rect 13461 3009 13495 3043
rect 15301 3009 15335 3043
rect 16681 3009 16715 3043
rect 16865 3009 16899 3043
rect 17049 3009 17083 3043
rect 17877 3009 17911 3043
rect 19717 3009 19751 3043
rect 19901 3009 19935 3043
rect 20085 3009 20119 3043
rect 20729 3009 20763 3043
rect 21005 3009 21039 3043
rect 21097 3009 21131 3043
rect 22293 3009 22327 3043
rect 23121 3009 23155 3043
rect 23581 3009 23615 3043
rect 23765 3009 23799 3043
rect 23949 3009 23983 3043
rect 25053 3009 25087 3043
rect 25320 3009 25354 3043
rect 27353 3009 27387 3043
rect 29653 3009 29687 3043
rect 29920 3009 29954 3043
rect 32137 3009 32171 3043
rect 32404 3009 32438 3043
rect 33977 3009 34011 3043
rect 35817 3009 35851 3043
rect 36737 3009 36771 3043
rect 37289 3009 37323 3043
rect 10609 2941 10643 2975
rect 22477 2941 22511 2975
rect 37565 2941 37599 2975
rect 3249 2873 3283 2907
rect 12081 2873 12115 2907
rect 14841 2873 14875 2907
rect 1593 2805 1627 2839
rect 2329 2805 2363 2839
rect 3065 2805 3099 2839
rect 5641 2805 5675 2839
rect 17233 2805 17267 2839
rect 20269 2805 20303 2839
rect 21281 2805 21315 2839
rect 24133 2805 24167 2839
rect 31033 2805 31067 2839
rect 33517 2805 33551 2839
rect 35357 2805 35391 2839
rect 36001 2805 36035 2839
rect 2651 2601 2685 2635
rect 14841 2601 14875 2635
rect 17049 2601 17083 2635
rect 19625 2601 19659 2635
rect 21005 2601 21039 2635
rect 23673 2601 23707 2635
rect 24869 2601 24903 2635
rect 28457 2601 28491 2635
rect 30205 2601 30239 2635
rect 31401 2601 31435 2635
rect 32505 2601 32539 2635
rect 22753 2533 22787 2567
rect 25881 2533 25915 2567
rect 34897 2533 34931 2567
rect 1961 2465 1995 2499
rect 2421 2465 2455 2499
rect 5273 2465 5307 2499
rect 16681 2465 16715 2499
rect 19257 2465 19291 2499
rect 20637 2465 20671 2499
rect 23305 2465 23339 2499
rect 24501 2465 24535 2499
rect 32137 2465 32171 2499
rect 37565 2465 37599 2499
rect 3985 2397 4019 2431
rect 4997 2397 5031 2431
rect 6929 2397 6963 2431
rect 7849 2397 7883 2431
rect 8953 2397 8987 2431
rect 9873 2397 9907 2431
rect 10793 2397 10827 2431
rect 11529 2397 11563 2431
rect 12265 2397 12299 2431
rect 13185 2397 13219 2431
rect 14289 2397 14323 2431
rect 14473 2397 14507 2431
rect 14657 2397 14691 2431
rect 15853 2397 15887 2431
rect 16865 2397 16899 2431
rect 17693 2397 17727 2431
rect 18429 2397 18463 2431
rect 19441 2397 19475 2431
rect 20821 2397 20855 2431
rect 21833 2397 21867 2431
rect 22569 2397 22603 2431
rect 23489 2397 23523 2431
rect 24685 2397 24719 2431
rect 25329 2397 25363 2431
rect 25697 2397 25731 2431
rect 26991 2397 27025 2431
rect 27905 2397 27939 2431
rect 28089 2397 28123 2431
rect 28273 2397 28307 2431
rect 29653 2397 29687 2431
rect 30021 2397 30055 2431
rect 30665 2397 30699 2431
rect 31585 2397 31619 2431
rect 32321 2397 32355 2431
rect 32965 2397 32999 2431
rect 33701 2397 33735 2431
rect 34713 2397 34747 2431
rect 35909 2397 35943 2431
rect 36185 2397 36219 2431
rect 37289 2397 37323 2431
rect 1777 2329 1811 2363
rect 14565 2329 14599 2363
rect 25513 2329 25547 2363
rect 25605 2329 25639 2363
rect 28181 2329 28215 2363
rect 29837 2329 29871 2363
rect 29929 2329 29963 2363
rect 4169 2261 4203 2295
rect 7113 2261 7147 2295
rect 7665 2261 7699 2295
rect 9137 2261 9171 2295
rect 10057 2261 10091 2295
rect 10609 2261 10643 2295
rect 11713 2261 11747 2295
rect 12449 2261 12483 2295
rect 13369 2261 13403 2295
rect 16037 2261 16071 2295
rect 17877 2261 17911 2295
rect 18613 2261 18647 2295
rect 22017 2261 22051 2295
rect 27169 2261 27203 2295
rect 30849 2261 30883 2295
rect 33149 2261 33183 2295
rect 33885 2261 33919 2295
<< metal1 >>
rect 2130 48152 2136 48204
rect 2188 48192 2194 48204
rect 13998 48192 14004 48204
rect 2188 48164 14004 48192
rect 2188 48152 2194 48164
rect 13998 48152 14004 48164
rect 14056 48152 14062 48204
rect 3602 48084 3608 48136
rect 3660 48124 3666 48136
rect 13170 48124 13176 48136
rect 3660 48096 13176 48124
rect 3660 48084 3666 48096
rect 13170 48084 13176 48096
rect 13228 48084 13234 48136
rect 3786 48016 3792 48068
rect 3844 48056 3850 48068
rect 15102 48056 15108 48068
rect 3844 48028 15108 48056
rect 3844 48016 3850 48028
rect 15102 48016 15108 48028
rect 15160 48016 15166 48068
rect 12986 47948 12992 48000
rect 13044 47988 13050 48000
rect 22462 47988 22468 48000
rect 13044 47960 22468 47988
rect 13044 47948 13050 47960
rect 22462 47948 22468 47960
rect 22520 47948 22526 48000
rect 10410 47880 10416 47932
rect 10468 47920 10474 47932
rect 20254 47920 20260 47932
rect 10468 47892 20260 47920
rect 10468 47880 10474 47892
rect 20254 47880 20260 47892
rect 20312 47880 20318 47932
rect 6362 47744 6368 47796
rect 6420 47784 6426 47796
rect 17494 47784 17500 47796
rect 6420 47756 17500 47784
rect 6420 47744 6426 47756
rect 17494 47744 17500 47756
rect 17552 47744 17558 47796
rect 5074 47676 5080 47728
rect 5132 47716 5138 47728
rect 16298 47716 16304 47728
rect 5132 47688 16304 47716
rect 5132 47676 5138 47688
rect 16298 47676 16304 47688
rect 16356 47676 16362 47728
rect 1394 47608 1400 47660
rect 1452 47648 1458 47660
rect 12066 47648 12072 47660
rect 1452 47620 12072 47648
rect 1452 47608 1458 47620
rect 12066 47608 12072 47620
rect 12124 47608 12130 47660
rect 12710 47608 12716 47660
rect 12768 47648 12774 47660
rect 27522 47648 27528 47660
rect 12768 47620 27528 47648
rect 12768 47608 12774 47620
rect 27522 47608 27528 47620
rect 27580 47608 27586 47660
rect 8938 47540 8944 47592
rect 8996 47580 9002 47592
rect 19978 47580 19984 47592
rect 8996 47552 19984 47580
rect 8996 47540 9002 47552
rect 19978 47540 19984 47552
rect 20036 47540 20042 47592
rect 5258 47472 5264 47524
rect 5316 47512 5322 47524
rect 17126 47512 17132 47524
rect 5316 47484 17132 47512
rect 5316 47472 5322 47484
rect 17126 47472 17132 47484
rect 17184 47472 17190 47524
rect 7098 47404 7104 47456
rect 7156 47444 7162 47456
rect 13906 47444 13912 47456
rect 7156 47416 13912 47444
rect 7156 47404 7162 47416
rect 13906 47404 13912 47416
rect 13964 47404 13970 47456
rect 20530 47404 20536 47456
rect 20588 47444 20594 47456
rect 30742 47444 30748 47456
rect 20588 47416 30748 47444
rect 20588 47404 20594 47416
rect 30742 47404 30748 47416
rect 30800 47404 30806 47456
rect 1104 47354 38824 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 38824 47354
rect 1104 47280 38824 47302
rect 382 47200 388 47252
rect 440 47240 446 47252
rect 1581 47243 1639 47249
rect 1581 47240 1593 47243
rect 440 47212 1593 47240
rect 440 47200 446 47212
rect 1581 47209 1593 47212
rect 1627 47209 1639 47243
rect 1581 47203 1639 47209
rect 2314 47200 2320 47252
rect 2372 47240 2378 47252
rect 3053 47243 3111 47249
rect 3053 47240 3065 47243
rect 2372 47212 3065 47240
rect 2372 47200 2378 47212
rect 3053 47209 3065 47212
rect 3099 47209 3111 47243
rect 3053 47203 3111 47209
rect 4614 47200 4620 47252
rect 4672 47240 4678 47252
rect 5445 47243 5503 47249
rect 5445 47240 5457 47243
rect 4672 47212 5457 47240
rect 4672 47200 4678 47212
rect 5445 47209 5457 47212
rect 5491 47209 5503 47243
rect 6546 47240 6552 47252
rect 6507 47212 6552 47240
rect 5445 47203 5503 47209
rect 6546 47200 6552 47212
rect 6604 47200 6610 47252
rect 7282 47240 7288 47252
rect 7243 47212 7288 47240
rect 7282 47200 7288 47212
rect 7340 47200 7346 47252
rect 8110 47240 8116 47252
rect 8071 47212 8116 47240
rect 8110 47200 8116 47212
rect 8168 47200 8174 47252
rect 8662 47200 8668 47252
rect 8720 47240 8726 47252
rect 9125 47243 9183 47249
rect 9125 47240 9137 47243
rect 8720 47212 9137 47240
rect 8720 47200 8726 47212
rect 9125 47209 9137 47212
rect 9171 47209 9183 47243
rect 9125 47203 9183 47209
rect 9674 47200 9680 47252
rect 9732 47240 9738 47252
rect 9861 47243 9919 47249
rect 9861 47240 9873 47243
rect 9732 47212 9873 47240
rect 9732 47200 9738 47212
rect 9861 47209 9873 47212
rect 9907 47209 9919 47243
rect 10594 47240 10600 47252
rect 10555 47212 10600 47240
rect 9861 47203 9919 47209
rect 10594 47200 10600 47212
rect 10652 47200 10658 47252
rect 11146 47200 11152 47252
rect 11204 47240 11210 47252
rect 11701 47243 11759 47249
rect 11701 47240 11713 47243
rect 11204 47212 11713 47240
rect 11204 47200 11210 47212
rect 11701 47209 11713 47212
rect 11747 47209 11759 47243
rect 11701 47203 11759 47209
rect 12434 47200 12440 47252
rect 12492 47240 12498 47252
rect 12492 47212 12537 47240
rect 12492 47200 12498 47212
rect 12802 47200 12808 47252
rect 12860 47240 12866 47252
rect 13173 47243 13231 47249
rect 13173 47240 13185 47243
rect 12860 47212 13185 47240
rect 12860 47200 12866 47212
rect 13173 47209 13185 47212
rect 13219 47209 13231 47243
rect 13173 47203 13231 47209
rect 13814 47200 13820 47252
rect 13872 47240 13878 47252
rect 14277 47243 14335 47249
rect 14277 47240 14289 47243
rect 13872 47212 14289 47240
rect 13872 47200 13878 47212
rect 14277 47209 14289 47212
rect 14323 47209 14335 47243
rect 14277 47203 14335 47209
rect 14550 47200 14556 47252
rect 14608 47240 14614 47252
rect 15013 47243 15071 47249
rect 15013 47240 15025 47243
rect 14608 47212 15025 47240
rect 14608 47200 14614 47212
rect 15013 47209 15025 47212
rect 15059 47209 15071 47243
rect 15013 47203 15071 47209
rect 15378 47200 15384 47252
rect 15436 47240 15442 47252
rect 15749 47243 15807 47249
rect 15749 47240 15761 47243
rect 15436 47212 15761 47240
rect 15436 47200 15442 47212
rect 15749 47209 15761 47212
rect 15795 47209 15807 47243
rect 15749 47203 15807 47209
rect 17034 47200 17040 47252
rect 17092 47240 17098 47252
rect 17589 47243 17647 47249
rect 17589 47240 17601 47243
rect 17092 47212 17601 47240
rect 17092 47200 17098 47212
rect 17589 47209 17601 47212
rect 17635 47209 17647 47243
rect 17589 47203 17647 47209
rect 17954 47200 17960 47252
rect 18012 47240 18018 47252
rect 18325 47243 18383 47249
rect 18325 47240 18337 47243
rect 18012 47212 18337 47240
rect 18012 47200 18018 47212
rect 18325 47209 18337 47212
rect 18371 47209 18383 47243
rect 18325 47203 18383 47209
rect 19518 47200 19524 47252
rect 19576 47240 19582 47252
rect 20165 47243 20223 47249
rect 20165 47240 20177 47243
rect 19576 47212 20177 47240
rect 19576 47200 19582 47212
rect 20165 47209 20177 47212
rect 20211 47209 20223 47243
rect 20165 47203 20223 47209
rect 20714 47200 20720 47252
rect 20772 47240 20778 47252
rect 20901 47243 20959 47249
rect 20901 47240 20913 47243
rect 20772 47212 20913 47240
rect 20772 47200 20778 47212
rect 20901 47209 20913 47212
rect 20947 47209 20959 47243
rect 20901 47203 20959 47209
rect 22094 47200 22100 47252
rect 22152 47240 22158 47252
rect 22281 47243 22339 47249
rect 22281 47240 22293 47243
rect 22152 47212 22293 47240
rect 22152 47200 22158 47212
rect 22281 47209 22293 47212
rect 22327 47209 22339 47243
rect 23106 47240 23112 47252
rect 23067 47212 23112 47240
rect 22281 47203 22339 47209
rect 23106 47200 23112 47212
rect 23164 47200 23170 47252
rect 23658 47200 23664 47252
rect 23716 47240 23722 47252
rect 24581 47243 24639 47249
rect 24581 47240 24593 47243
rect 23716 47212 24593 47240
rect 23716 47200 23722 47212
rect 24581 47209 24593 47212
rect 24627 47209 24639 47243
rect 24581 47203 24639 47209
rect 25314 47200 25320 47252
rect 25372 47240 25378 47252
rect 26053 47243 26111 47249
rect 26053 47240 26065 47243
rect 25372 47212 26065 47240
rect 25372 47200 25378 47212
rect 26053 47209 26065 47212
rect 26099 47209 26111 47243
rect 27522 47240 27528 47252
rect 27483 47212 27528 47240
rect 26053 47203 26111 47209
rect 27522 47200 27528 47212
rect 27580 47200 27586 47252
rect 30742 47200 30748 47252
rect 30800 47240 30806 47252
rect 35345 47243 35403 47249
rect 35345 47240 35357 47243
rect 30800 47212 35357 47240
rect 30800 47200 30806 47212
rect 35345 47209 35357 47212
rect 35391 47209 35403 47243
rect 35345 47203 35403 47209
rect 3970 47132 3976 47184
rect 4028 47172 4034 47184
rect 4709 47175 4767 47181
rect 4709 47172 4721 47175
rect 4028 47144 4721 47172
rect 4028 47132 4034 47144
rect 4709 47141 4721 47144
rect 4755 47141 4767 47175
rect 21082 47172 21088 47184
rect 4709 47135 4767 47141
rect 9692 47144 21088 47172
rect 1394 47036 1400 47048
rect 1355 47008 1400 47036
rect 1394 46996 1400 47008
rect 1452 46996 1458 47048
rect 2130 47036 2136 47048
rect 2091 47008 2136 47036
rect 2130 46996 2136 47008
rect 2188 46996 2194 47048
rect 2869 47039 2927 47045
rect 2869 47005 2881 47039
rect 2915 47036 2927 47039
rect 3602 47036 3608 47048
rect 2915 47008 3608 47036
rect 2915 47005 2927 47008
rect 2869 46999 2927 47005
rect 3602 46996 3608 47008
rect 3660 46996 3666 47048
rect 3786 47036 3792 47048
rect 3747 47008 3792 47036
rect 3786 46996 3792 47008
rect 3844 46996 3850 47048
rect 4525 47039 4583 47045
rect 4525 47005 4537 47039
rect 4571 47036 4583 47039
rect 5074 47036 5080 47048
rect 4571 47008 5080 47036
rect 4571 47005 4583 47008
rect 4525 46999 4583 47005
rect 5074 46996 5080 47008
rect 5132 46996 5138 47048
rect 5258 47036 5264 47048
rect 5219 47008 5264 47036
rect 5258 46996 5264 47008
rect 5316 46996 5322 47048
rect 6362 47036 6368 47048
rect 6323 47008 6368 47036
rect 6362 46996 6368 47008
rect 6420 46996 6426 47048
rect 7098 47036 7104 47048
rect 7059 47008 7104 47036
rect 7098 46996 7104 47008
rect 7156 46996 7162 47048
rect 7929 47039 7987 47045
rect 7929 47005 7941 47039
rect 7975 47005 7987 47039
rect 8938 47036 8944 47048
rect 8899 47008 8944 47036
rect 7929 46999 7987 47005
rect 1210 46928 1216 46980
rect 1268 46968 1274 46980
rect 1268 46940 2360 46968
rect 1268 46928 1274 46940
rect 2332 46909 2360 46940
rect 2958 46928 2964 46980
rect 3016 46968 3022 46980
rect 7944 46968 7972 46999
rect 8938 46996 8944 47008
rect 8996 46996 9002 47048
rect 9692 47045 9720 47144
rect 21082 47132 21088 47144
rect 21140 47132 21146 47184
rect 31018 47132 31024 47184
rect 31076 47172 31082 47184
rect 31297 47175 31355 47181
rect 31297 47172 31309 47175
rect 31076 47144 31309 47172
rect 31076 47132 31082 47144
rect 31297 47141 31309 47144
rect 31343 47141 31355 47175
rect 31297 47135 31355 47141
rect 12268 47076 17264 47104
rect 9677 47039 9735 47045
rect 9677 47005 9689 47039
rect 9723 47005 9735 47039
rect 10410 47036 10416 47048
rect 10371 47008 10416 47036
rect 9677 46999 9735 47005
rect 10410 46996 10416 47008
rect 10468 46996 10474 47048
rect 11514 47036 11520 47048
rect 11475 47008 11520 47036
rect 11514 46996 11520 47008
rect 11572 46996 11578 47048
rect 12268 47045 12296 47076
rect 12253 47039 12311 47045
rect 12253 47005 12265 47039
rect 12299 47005 12311 47039
rect 12986 47036 12992 47048
rect 12947 47008 12992 47036
rect 12253 46999 12311 47005
rect 12986 46996 12992 47008
rect 13044 46996 13050 47048
rect 13262 46996 13268 47048
rect 13320 47036 13326 47048
rect 14093 47039 14151 47045
rect 14093 47036 14105 47039
rect 13320 47008 14105 47036
rect 13320 46996 13326 47008
rect 14093 47005 14105 47008
rect 14139 47005 14151 47039
rect 14826 47036 14832 47048
rect 14787 47008 14832 47036
rect 14093 46999 14151 47005
rect 14826 46996 14832 47008
rect 14884 46996 14890 47048
rect 15562 47036 15568 47048
rect 15523 47008 15568 47036
rect 15562 46996 15568 47008
rect 15620 46996 15626 47048
rect 16574 46996 16580 47048
rect 16632 47036 16638 47048
rect 16669 47039 16727 47045
rect 16669 47036 16681 47039
rect 16632 47008 16681 47036
rect 16632 46996 16638 47008
rect 16669 47005 16681 47008
rect 16715 47005 16727 47039
rect 16669 46999 16727 47005
rect 17236 46968 17264 47076
rect 28166 47064 28172 47116
rect 28224 47104 28230 47116
rect 28353 47107 28411 47113
rect 28353 47104 28365 47107
rect 28224 47076 28365 47104
rect 28224 47064 28230 47076
rect 28353 47073 28365 47076
rect 28399 47073 28411 47107
rect 28353 47067 28411 47073
rect 28994 47064 29000 47116
rect 29052 47104 29058 47116
rect 29549 47107 29607 47113
rect 29549 47104 29561 47107
rect 29052 47076 29561 47104
rect 29052 47064 29058 47076
rect 29549 47073 29561 47076
rect 29595 47073 29607 47107
rect 29549 47067 29607 47073
rect 35894 47064 35900 47116
rect 35952 47104 35958 47116
rect 37277 47107 37335 47113
rect 35952 47076 35997 47104
rect 35952 47064 35958 47076
rect 37277 47073 37289 47107
rect 37323 47104 37335 47107
rect 37826 47104 37832 47116
rect 37323 47076 37832 47104
rect 37323 47073 37335 47076
rect 37277 47067 37335 47073
rect 37826 47064 37832 47076
rect 37884 47064 37890 47116
rect 17402 47036 17408 47048
rect 17363 47008 17408 47036
rect 17402 46996 17408 47008
rect 17460 46996 17466 47048
rect 18138 47036 18144 47048
rect 18099 47008 18144 47036
rect 18138 46996 18144 47008
rect 18196 46996 18202 47048
rect 18230 46996 18236 47048
rect 18288 47036 18294 47048
rect 19245 47039 19303 47045
rect 19245 47036 19257 47039
rect 18288 47008 19257 47036
rect 18288 46996 18294 47008
rect 19245 47005 19257 47008
rect 19291 47005 19303 47039
rect 19245 46999 19303 47005
rect 19334 46996 19340 47048
rect 19392 47036 19398 47048
rect 19981 47039 20039 47045
rect 19981 47036 19993 47039
rect 19392 47008 19993 47036
rect 19392 46996 19398 47008
rect 19981 47005 19993 47008
rect 20027 47005 20039 47039
rect 20714 47036 20720 47048
rect 20675 47008 20720 47036
rect 19981 46999 20039 47005
rect 20714 46996 20720 47008
rect 20772 46996 20778 47048
rect 22094 47036 22100 47048
rect 22055 47008 22100 47036
rect 22094 46996 22100 47008
rect 22152 46996 22158 47048
rect 22922 47036 22928 47048
rect 22883 47008 22928 47036
rect 22922 46996 22928 47008
rect 22980 46996 22986 47048
rect 24394 47036 24400 47048
rect 24355 47008 24400 47036
rect 24394 46996 24400 47008
rect 24452 46996 24458 47048
rect 25133 47039 25191 47045
rect 25133 47036 25145 47039
rect 24504 47008 25145 47036
rect 23382 46968 23388 46980
rect 3016 46940 4016 46968
rect 7944 46940 17172 46968
rect 17236 46940 23388 46968
rect 3016 46928 3022 46940
rect 3988 46909 4016 46940
rect 2317 46903 2375 46909
rect 2317 46869 2329 46903
rect 2363 46869 2375 46903
rect 2317 46863 2375 46869
rect 3973 46903 4031 46909
rect 3973 46869 3985 46903
rect 4019 46869 4031 46903
rect 3973 46863 4031 46869
rect 16206 46860 16212 46912
rect 16264 46900 16270 46912
rect 16853 46903 16911 46909
rect 16853 46900 16865 46903
rect 16264 46872 16865 46900
rect 16264 46860 16270 46872
rect 16853 46869 16865 46872
rect 16899 46869 16911 46903
rect 17144 46900 17172 46940
rect 23382 46928 23388 46940
rect 23440 46928 23446 46980
rect 23934 46928 23940 46980
rect 23992 46968 23998 46980
rect 24504 46968 24532 47008
rect 25133 47005 25145 47008
rect 25179 47005 25191 47039
rect 25133 46999 25191 47005
rect 25869 47039 25927 47045
rect 25869 47005 25881 47039
rect 25915 47005 25927 47039
rect 25869 46999 25927 47005
rect 23992 46940 24532 46968
rect 23992 46928 23998 46940
rect 24578 46928 24584 46980
rect 24636 46968 24642 46980
rect 25884 46968 25912 46999
rect 27062 46996 27068 47048
rect 27120 47036 27126 47048
rect 27433 47039 27491 47045
rect 27433 47036 27445 47039
rect 27120 47008 27445 47036
rect 27120 46996 27126 47008
rect 27433 47005 27445 47008
rect 27479 47005 27491 47039
rect 29822 47036 29828 47048
rect 29783 47008 29828 47036
rect 27433 46999 27491 47005
rect 29822 46996 29828 47008
rect 29880 46996 29886 47048
rect 31478 47036 31484 47048
rect 31439 47008 31484 47036
rect 31478 46996 31484 47008
rect 31536 46996 31542 47048
rect 32125 47039 32183 47045
rect 32125 47036 32137 47039
rect 31772 47008 32137 47036
rect 24636 46940 25912 46968
rect 24636 46928 24642 46940
rect 27890 46928 27896 46980
rect 27948 46968 27954 46980
rect 28169 46971 28227 46977
rect 28169 46968 28181 46971
rect 27948 46940 28181 46968
rect 27948 46928 27954 46940
rect 28169 46937 28181 46940
rect 28215 46937 28227 46971
rect 28169 46931 28227 46937
rect 18046 46900 18052 46912
rect 17144 46872 18052 46900
rect 16853 46863 16911 46869
rect 18046 46860 18052 46872
rect 18104 46860 18110 46912
rect 18690 46860 18696 46912
rect 18748 46900 18754 46912
rect 19429 46903 19487 46909
rect 19429 46900 19441 46903
rect 18748 46872 19441 46900
rect 18748 46860 18754 46872
rect 19429 46869 19441 46872
rect 19475 46869 19487 46903
rect 19429 46863 19487 46869
rect 24486 46860 24492 46912
rect 24544 46900 24550 46912
rect 25317 46903 25375 46909
rect 25317 46900 25329 46903
rect 24544 46872 25329 46900
rect 24544 46860 24550 46872
rect 25317 46869 25329 46872
rect 25363 46869 25375 46903
rect 25317 46863 25375 46869
rect 30374 46860 30380 46912
rect 30432 46900 30438 46912
rect 31772 46900 31800 47008
rect 32125 47005 32137 47008
rect 32171 47005 32183 47039
rect 32398 47036 32404 47048
rect 32359 47008 32404 47036
rect 32125 46999 32183 47005
rect 32398 46996 32404 47008
rect 32456 46996 32462 47048
rect 33870 47036 33876 47048
rect 33831 47008 33876 47036
rect 33870 46996 33876 47008
rect 33928 46996 33934 47048
rect 35253 47039 35311 47045
rect 35253 47005 35265 47039
rect 35299 47036 35311 47039
rect 35342 47036 35348 47048
rect 35299 47008 35348 47036
rect 35299 47005 35311 47008
rect 35253 46999 35311 47005
rect 35342 46996 35348 47008
rect 35400 46996 35406 47048
rect 36170 47036 36176 47048
rect 36131 47008 36176 47036
rect 36170 46996 36176 47008
rect 36228 46996 36234 47048
rect 37550 47036 37556 47048
rect 37511 47008 37556 47036
rect 37550 46996 37556 47008
rect 37608 46996 37614 47048
rect 34054 46968 34060 46980
rect 34015 46940 34060 46968
rect 34054 46928 34060 46940
rect 34112 46928 34118 46980
rect 30432 46872 31800 46900
rect 30432 46860 30438 46872
rect 1104 46810 38824 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 38824 46810
rect 1104 46736 38824 46758
rect 5350 46656 5356 46708
rect 5408 46696 5414 46708
rect 5629 46699 5687 46705
rect 5629 46696 5641 46699
rect 5408 46668 5641 46696
rect 5408 46656 5414 46668
rect 5629 46665 5641 46668
rect 5675 46665 5687 46699
rect 5629 46659 5687 46665
rect 12161 46699 12219 46705
rect 12161 46665 12173 46699
rect 12207 46696 12219 46699
rect 13262 46696 13268 46708
rect 12207 46668 13268 46696
rect 12207 46665 12219 46668
rect 12161 46659 12219 46665
rect 13262 46656 13268 46668
rect 13320 46656 13326 46708
rect 14277 46699 14335 46705
rect 14277 46665 14289 46699
rect 14323 46696 14335 46699
rect 15562 46696 15568 46708
rect 14323 46668 15568 46696
rect 14323 46665 14335 46668
rect 14277 46659 14335 46665
rect 15562 46656 15568 46668
rect 15620 46656 15626 46708
rect 15933 46699 15991 46705
rect 15933 46665 15945 46699
rect 15979 46696 15991 46699
rect 17402 46696 17408 46708
rect 15979 46668 17408 46696
rect 15979 46665 15991 46668
rect 15933 46659 15991 46665
rect 17402 46656 17408 46668
rect 17460 46656 17466 46708
rect 17681 46699 17739 46705
rect 17681 46665 17693 46699
rect 17727 46696 17739 46699
rect 18230 46696 18236 46708
rect 17727 46668 18236 46696
rect 17727 46665 17739 46668
rect 17681 46659 17739 46665
rect 18230 46656 18236 46668
rect 18288 46656 18294 46708
rect 18509 46699 18567 46705
rect 18509 46665 18521 46699
rect 18555 46696 18567 46699
rect 19334 46696 19340 46708
rect 18555 46668 19340 46696
rect 18555 46665 18567 46668
rect 18509 46659 18567 46665
rect 19334 46656 19340 46668
rect 19392 46656 19398 46708
rect 19521 46699 19579 46705
rect 19521 46665 19533 46699
rect 19567 46696 19579 46699
rect 20714 46696 20720 46708
rect 19567 46668 20720 46696
rect 19567 46665 19579 46668
rect 19521 46659 19579 46665
rect 20714 46656 20720 46668
rect 20772 46656 20778 46708
rect 20993 46699 21051 46705
rect 20993 46665 21005 46699
rect 21039 46696 21051 46699
rect 22094 46696 22100 46708
rect 21039 46668 22100 46696
rect 21039 46665 21051 46668
rect 20993 46659 21051 46665
rect 22094 46656 22100 46668
rect 22152 46656 22158 46708
rect 23845 46699 23903 46705
rect 23845 46665 23857 46699
rect 23891 46665 23903 46699
rect 23845 46659 23903 46665
rect 13817 46631 13875 46637
rect 13817 46628 13829 46631
rect 13004 46600 13829 46628
rect 5442 46560 5448 46572
rect 5403 46532 5448 46560
rect 5442 46520 5448 46532
rect 5500 46520 5506 46572
rect 12250 46520 12256 46572
rect 12308 46560 12314 46572
rect 13004 46569 13032 46600
rect 13817 46597 13829 46600
rect 13863 46597 13875 46631
rect 17037 46631 17095 46637
rect 17037 46628 17049 46631
rect 13817 46591 13875 46597
rect 15488 46600 17049 46628
rect 12345 46563 12403 46569
rect 12345 46560 12357 46563
rect 12308 46532 12357 46560
rect 12308 46520 12314 46532
rect 12345 46529 12357 46532
rect 12391 46529 12403 46563
rect 12345 46523 12403 46529
rect 12989 46563 13047 46569
rect 12989 46529 13001 46563
rect 13035 46529 13047 46563
rect 12989 46523 13047 46529
rect 13633 46563 13691 46569
rect 13633 46529 13645 46563
rect 13679 46560 13691 46563
rect 13998 46560 14004 46572
rect 13679 46532 14004 46560
rect 13679 46529 13691 46532
rect 13633 46523 13691 46529
rect 13998 46520 14004 46532
rect 14056 46520 14062 46572
rect 14458 46560 14464 46572
rect 14419 46532 14464 46560
rect 14458 46520 14464 46532
rect 14516 46520 14522 46572
rect 15488 46569 15516 46600
rect 17037 46597 17049 46600
rect 17083 46597 17095 46631
rect 21358 46628 21364 46640
rect 17037 46591 17095 46597
rect 17328 46600 21364 46628
rect 15473 46563 15531 46569
rect 15473 46529 15485 46563
rect 15519 46529 15531 46563
rect 15473 46523 15531 46529
rect 16117 46563 16175 46569
rect 16117 46529 16129 46563
rect 16163 46560 16175 46563
rect 16482 46560 16488 46572
rect 16163 46532 16488 46560
rect 16163 46529 16175 46532
rect 16117 46523 16175 46529
rect 16482 46520 16488 46532
rect 16540 46520 16546 46572
rect 17328 46569 17356 46600
rect 21358 46588 21364 46600
rect 21416 46588 21422 46640
rect 23860 46628 23888 46659
rect 26142 46656 26148 46708
rect 26200 46696 26206 46708
rect 27157 46699 27215 46705
rect 27157 46696 27169 46699
rect 26200 46668 27169 46696
rect 26200 46656 26206 46668
rect 27157 46665 27169 46668
rect 27203 46665 27215 46699
rect 27157 46659 27215 46665
rect 34698 46628 34704 46640
rect 23860 46600 26234 46628
rect 34659 46600 34704 46628
rect 16853 46563 16911 46569
rect 16853 46560 16865 46563
rect 16592 46532 16865 46560
rect 11698 46452 11704 46504
rect 11756 46492 11762 46504
rect 13449 46495 13507 46501
rect 13449 46492 13461 46495
rect 11756 46464 13461 46492
rect 11756 46452 11762 46464
rect 13449 46461 13461 46464
rect 13495 46461 13507 46495
rect 13449 46455 13507 46461
rect 15102 46452 15108 46504
rect 15160 46492 15166 46504
rect 16592 46492 16620 46532
rect 16853 46529 16865 46532
rect 16899 46560 16911 46563
rect 17313 46563 17371 46569
rect 17313 46560 17325 46563
rect 16899 46532 17325 46560
rect 16899 46529 16911 46532
rect 16853 46523 16911 46529
rect 17313 46529 17325 46532
rect 17359 46529 17371 46563
rect 17862 46560 17868 46572
rect 17823 46532 17868 46560
rect 17313 46523 17371 46529
rect 17862 46520 17868 46532
rect 17920 46520 17926 46572
rect 18690 46560 18696 46572
rect 18651 46532 18696 46560
rect 18690 46520 18696 46532
rect 18748 46520 18754 46572
rect 19705 46563 19763 46569
rect 19705 46560 19717 46563
rect 18800 46532 19717 46560
rect 15160 46464 16620 46492
rect 16669 46495 16727 46501
rect 15160 46452 15166 46464
rect 16669 46461 16681 46495
rect 16715 46492 16727 46495
rect 17770 46492 17776 46504
rect 16715 46464 17776 46492
rect 16715 46461 16727 46464
rect 16669 46455 16727 46461
rect 17770 46452 17776 46464
rect 17828 46452 17834 46504
rect 12805 46427 12863 46433
rect 12805 46393 12817 46427
rect 12851 46424 12863 46427
rect 14826 46424 14832 46436
rect 12851 46396 14832 46424
rect 12851 46393 12863 46396
rect 12805 46387 12863 46393
rect 14826 46384 14832 46396
rect 14884 46384 14890 46436
rect 15289 46427 15347 46433
rect 15289 46393 15301 46427
rect 15335 46424 15347 46427
rect 16574 46424 16580 46436
rect 15335 46396 16580 46424
rect 15335 46393 15347 46396
rect 15289 46387 15347 46393
rect 16574 46384 16580 46396
rect 16632 46384 16638 46436
rect 18800 46424 18828 46532
rect 19705 46529 19717 46532
rect 19751 46529 19763 46563
rect 21174 46560 21180 46572
rect 21135 46532 21180 46560
rect 19705 46523 19763 46529
rect 21174 46520 21180 46532
rect 21232 46520 21238 46572
rect 21821 46563 21879 46569
rect 21821 46529 21833 46563
rect 21867 46529 21879 46563
rect 24026 46560 24032 46572
rect 23987 46532 24032 46560
rect 21821 46523 21879 46529
rect 19334 46452 19340 46504
rect 19392 46492 19398 46504
rect 21836 46492 21864 46523
rect 24026 46520 24032 46532
rect 24084 46520 24090 46572
rect 26206 46560 26234 46600
rect 34698 46588 34704 46600
rect 34756 46588 34762 46640
rect 26973 46563 27031 46569
rect 26973 46560 26985 46563
rect 26206 46532 26985 46560
rect 26973 46529 26985 46532
rect 27019 46529 27031 46563
rect 29638 46560 29644 46572
rect 29599 46532 29644 46560
rect 26973 46523 27031 46529
rect 29638 46520 29644 46532
rect 29696 46520 29702 46572
rect 32306 46560 32312 46572
rect 32267 46532 32312 46560
rect 32306 46520 32312 46532
rect 32364 46520 32370 46572
rect 32858 46520 32864 46572
rect 32916 46560 32922 46572
rect 33137 46563 33195 46569
rect 33137 46560 33149 46563
rect 32916 46532 33149 46560
rect 32916 46520 32922 46532
rect 33137 46529 33149 46532
rect 33183 46529 33195 46563
rect 33137 46523 33195 46529
rect 37277 46563 37335 46569
rect 37277 46529 37289 46563
rect 37323 46560 37335 46563
rect 38654 46560 38660 46572
rect 37323 46532 38660 46560
rect 37323 46529 37335 46532
rect 37277 46523 37335 46529
rect 38654 46520 38660 46532
rect 38712 46520 38718 46572
rect 29914 46492 29920 46504
rect 19392 46464 21864 46492
rect 29875 46464 29920 46492
rect 19392 46452 19398 46464
rect 29914 46452 29920 46464
rect 29972 46452 29978 46504
rect 37458 46452 37464 46504
rect 37516 46492 37522 46504
rect 37553 46495 37611 46501
rect 37553 46492 37565 46495
rect 37516 46464 37565 46492
rect 37516 46452 37522 46464
rect 37553 46461 37565 46464
rect 37599 46461 37611 46495
rect 37553 46455 37611 46461
rect 16684 46396 18828 46424
rect 14918 46316 14924 46368
rect 14976 46356 14982 46368
rect 16684 46356 16712 46396
rect 21266 46384 21272 46436
rect 21324 46424 21330 46436
rect 22005 46427 22063 46433
rect 22005 46424 22017 46427
rect 21324 46396 22017 46424
rect 21324 46384 21330 46396
rect 22005 46393 22017 46396
rect 22051 46393 22063 46427
rect 22005 46387 22063 46393
rect 32122 46356 32128 46368
rect 14976 46328 16712 46356
rect 32083 46328 32128 46356
rect 14976 46316 14982 46328
rect 32122 46316 32128 46328
rect 32180 46316 32186 46368
rect 32950 46356 32956 46368
rect 32911 46328 32956 46356
rect 32950 46316 32956 46328
rect 33008 46316 33014 46368
rect 34790 46356 34796 46368
rect 34751 46328 34796 46356
rect 34790 46316 34796 46328
rect 34848 46316 34854 46368
rect 1104 46266 38824 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 38824 46266
rect 1104 46192 38824 46214
rect 5442 46112 5448 46164
rect 5500 46152 5506 46164
rect 12250 46152 12256 46164
rect 5500 46124 6914 46152
rect 12211 46124 12256 46152
rect 5500 46112 5506 46124
rect 6886 45880 6914 46124
rect 12250 46112 12256 46124
rect 12308 46112 12314 46164
rect 13449 46155 13507 46161
rect 13449 46121 13461 46155
rect 13495 46152 13507 46155
rect 14458 46152 14464 46164
rect 13495 46124 14464 46152
rect 13495 46121 13507 46124
rect 13449 46115 13507 46121
rect 14458 46112 14464 46124
rect 14516 46112 14522 46164
rect 14829 46155 14887 46161
rect 14829 46121 14841 46155
rect 14875 46152 14887 46155
rect 14918 46152 14924 46164
rect 14875 46124 14924 46152
rect 14875 46121 14887 46124
rect 14829 46115 14887 46121
rect 14918 46112 14924 46124
rect 14976 46112 14982 46164
rect 16482 46152 16488 46164
rect 16443 46124 16488 46152
rect 16482 46112 16488 46124
rect 16540 46112 16546 46164
rect 17773 46155 17831 46161
rect 17773 46121 17785 46155
rect 17819 46152 17831 46155
rect 18138 46152 18144 46164
rect 17819 46124 18144 46152
rect 17819 46121 17831 46124
rect 17773 46115 17831 46121
rect 18138 46112 18144 46124
rect 18196 46112 18202 46164
rect 22189 46155 22247 46161
rect 22189 46121 22201 46155
rect 22235 46152 22247 46155
rect 22922 46152 22928 46164
rect 22235 46124 22928 46152
rect 22235 46121 22247 46124
rect 22189 46115 22247 46121
rect 22922 46112 22928 46124
rect 22980 46112 22986 46164
rect 15657 46087 15715 46093
rect 15657 46053 15669 46087
rect 15703 46084 15715 46087
rect 17862 46084 17868 46096
rect 15703 46056 17868 46084
rect 15703 46053 15715 46056
rect 15657 46047 15715 46053
rect 17862 46044 17868 46056
rect 17920 46044 17926 46096
rect 10686 45976 10692 46028
rect 10744 46016 10750 46028
rect 13081 46019 13139 46025
rect 13081 46016 13093 46019
rect 10744 45988 13093 46016
rect 10744 45976 10750 45988
rect 13081 45985 13093 45988
rect 13127 45985 13139 46019
rect 13081 45979 13139 45985
rect 14090 45976 14096 46028
rect 14148 46016 14154 46028
rect 14148 45988 14780 46016
rect 14148 45976 14154 45988
rect 11974 45948 11980 45960
rect 11935 45920 11980 45948
rect 11974 45908 11980 45920
rect 12032 45908 12038 45960
rect 12066 45908 12072 45960
rect 12124 45948 12130 45960
rect 13262 45948 13268 45960
rect 12124 45920 12169 45948
rect 13223 45920 13268 45948
rect 12124 45908 12130 45920
rect 13262 45908 13268 45920
rect 13320 45908 13326 45960
rect 14458 45948 14464 45960
rect 14419 45920 14464 45948
rect 14458 45908 14464 45920
rect 14516 45908 14522 45960
rect 14645 45951 14703 45957
rect 14645 45917 14657 45951
rect 14691 45917 14703 45951
rect 14752 45948 14780 45988
rect 15102 45976 15108 46028
rect 15160 46016 15166 46028
rect 16117 46019 16175 46025
rect 16117 46016 16129 46019
rect 15160 45988 16129 46016
rect 15160 45976 15166 45988
rect 16117 45985 16129 45988
rect 16163 45985 16175 46019
rect 23290 46016 23296 46028
rect 16117 45979 16175 45985
rect 16960 45988 23296 46016
rect 15289 45951 15347 45957
rect 15289 45948 15301 45951
rect 14752 45920 15301 45948
rect 14645 45911 14703 45917
rect 15289 45917 15301 45920
rect 15335 45917 15347 45951
rect 15470 45948 15476 45960
rect 15431 45920 15476 45948
rect 15289 45911 15347 45917
rect 6886 45852 12434 45880
rect 12406 45812 12434 45852
rect 13906 45840 13912 45892
rect 13964 45880 13970 45892
rect 14660 45880 14688 45911
rect 15470 45908 15476 45920
rect 15528 45908 15534 45960
rect 16298 45948 16304 45960
rect 16211 45920 16304 45948
rect 16298 45908 16304 45920
rect 16356 45948 16362 45960
rect 16960 45948 16988 45988
rect 23290 45976 23296 45988
rect 23348 45976 23354 46028
rect 16356 45920 16988 45948
rect 17037 45951 17095 45957
rect 16356 45908 16362 45920
rect 17037 45917 17049 45951
rect 17083 45917 17095 45951
rect 17037 45911 17095 45917
rect 13964 45852 14688 45880
rect 17052 45880 17080 45911
rect 17126 45908 17132 45960
rect 17184 45948 17190 45960
rect 17313 45951 17371 45957
rect 17184 45920 17229 45948
rect 17184 45908 17190 45920
rect 17313 45917 17325 45951
rect 17359 45948 17371 45951
rect 17957 45951 18015 45957
rect 17957 45948 17969 45951
rect 17359 45920 17969 45948
rect 17359 45917 17371 45920
rect 17313 45911 17371 45917
rect 17957 45917 17969 45920
rect 18003 45917 18015 45951
rect 22370 45948 22376 45960
rect 22331 45920 22376 45948
rect 17957 45911 18015 45917
rect 22370 45908 22376 45920
rect 22428 45908 22434 45960
rect 37182 45948 37188 45960
rect 37143 45920 37188 45948
rect 37182 45908 37188 45920
rect 37240 45908 37246 45960
rect 37921 45951 37979 45957
rect 37921 45917 37933 45951
rect 37967 45948 37979 45951
rect 39482 45948 39488 45960
rect 37967 45920 39488 45948
rect 37967 45917 37979 45920
rect 37921 45911 37979 45917
rect 39482 45908 39488 45920
rect 39540 45908 39546 45960
rect 17218 45880 17224 45892
rect 17052 45852 17224 45880
rect 13964 45840 13970 45852
rect 17218 45840 17224 45852
rect 17276 45840 17282 45892
rect 15470 45812 15476 45824
rect 12406 45784 15476 45812
rect 15470 45772 15476 45784
rect 15528 45772 15534 45824
rect 37274 45812 37280 45824
rect 37235 45784 37280 45812
rect 37274 45772 37280 45784
rect 37332 45772 37338 45824
rect 38010 45812 38016 45824
rect 37971 45784 38016 45812
rect 38010 45772 38016 45784
rect 38068 45772 38074 45824
rect 1104 45722 38824 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 38824 45722
rect 1104 45648 38824 45670
rect 13262 45568 13268 45620
rect 13320 45608 13326 45620
rect 18138 45608 18144 45620
rect 13320 45580 18144 45608
rect 13320 45568 13326 45580
rect 18138 45568 18144 45580
rect 18196 45568 18202 45620
rect 23290 45608 23296 45620
rect 23251 45580 23296 45608
rect 23290 45568 23296 45580
rect 23348 45568 23354 45620
rect 17681 45543 17739 45549
rect 17681 45509 17693 45543
rect 17727 45540 17739 45543
rect 18690 45540 18696 45552
rect 17727 45512 18696 45540
rect 17727 45509 17739 45512
rect 17681 45503 17739 45509
rect 18690 45500 18696 45512
rect 18748 45500 18754 45552
rect 20165 45543 20223 45549
rect 20165 45509 20177 45543
rect 20211 45540 20223 45543
rect 21174 45540 21180 45552
rect 20211 45512 21180 45540
rect 20211 45509 20223 45512
rect 20165 45503 20223 45509
rect 21174 45500 21180 45512
rect 21232 45500 21238 45552
rect 21269 45543 21327 45549
rect 21269 45509 21281 45543
rect 21315 45540 21327 45543
rect 22370 45540 22376 45552
rect 21315 45512 22376 45540
rect 21315 45509 21327 45512
rect 21269 45503 21327 45509
rect 22370 45500 22376 45512
rect 22428 45500 22434 45552
rect 22649 45543 22707 45549
rect 22649 45509 22661 45543
rect 22695 45540 22707 45543
rect 24026 45540 24032 45552
rect 22695 45512 24032 45540
rect 22695 45509 22707 45512
rect 22649 45503 22707 45509
rect 24026 45500 24032 45512
rect 24084 45500 24090 45552
rect 12250 45432 12256 45484
rect 12308 45472 12314 45484
rect 13081 45475 13139 45481
rect 13081 45472 13093 45475
rect 12308 45444 13093 45472
rect 12308 45432 12314 45444
rect 13081 45441 13093 45444
rect 13127 45441 13139 45475
rect 13081 45435 13139 45441
rect 13817 45475 13875 45481
rect 13817 45441 13829 45475
rect 13863 45472 13875 45475
rect 13998 45472 14004 45484
rect 13863 45444 14004 45472
rect 13863 45441 13875 45444
rect 13817 45435 13875 45441
rect 13998 45432 14004 45444
rect 14056 45432 14062 45484
rect 17494 45472 17500 45484
rect 17455 45444 17500 45472
rect 17494 45432 17500 45444
rect 17552 45432 17558 45484
rect 18322 45432 18328 45484
rect 18380 45472 18386 45484
rect 19337 45475 19395 45481
rect 19337 45472 19349 45475
rect 18380 45444 19349 45472
rect 18380 45432 18386 45444
rect 19337 45441 19349 45444
rect 19383 45441 19395 45475
rect 19978 45472 19984 45484
rect 19939 45444 19984 45472
rect 19337 45435 19395 45441
rect 19978 45432 19984 45444
rect 20036 45432 20042 45484
rect 21082 45472 21088 45484
rect 21043 45444 21088 45472
rect 21082 45432 21088 45444
rect 21140 45432 21146 45484
rect 22462 45472 22468 45484
rect 22423 45444 22468 45472
rect 22462 45432 22468 45444
rect 22520 45432 22526 45484
rect 23201 45475 23259 45481
rect 23201 45441 23213 45475
rect 23247 45472 23259 45475
rect 24210 45472 24216 45484
rect 23247 45444 24216 45472
rect 23247 45441 23259 45444
rect 23201 45435 23259 45441
rect 24210 45432 24216 45444
rect 24268 45432 24274 45484
rect 29733 45475 29791 45481
rect 29733 45441 29745 45475
rect 29779 45472 29791 45475
rect 30374 45472 30380 45484
rect 29779 45444 30380 45472
rect 29779 45441 29791 45444
rect 29733 45435 29791 45441
rect 30374 45432 30380 45444
rect 30432 45432 30438 45484
rect 13538 45404 13544 45416
rect 13499 45376 13544 45404
rect 13538 45364 13544 45376
rect 13596 45364 13602 45416
rect 17310 45404 17316 45416
rect 17271 45376 17316 45404
rect 17310 45364 17316 45376
rect 17368 45364 17374 45416
rect 19797 45407 19855 45413
rect 19797 45373 19809 45407
rect 19843 45404 19855 45407
rect 20622 45404 20628 45416
rect 19843 45376 20628 45404
rect 19843 45373 19855 45376
rect 19797 45367 19855 45373
rect 20622 45364 20628 45376
rect 20680 45364 20686 45416
rect 20901 45407 20959 45413
rect 20901 45373 20913 45407
rect 20947 45404 20959 45407
rect 22281 45407 22339 45413
rect 20947 45376 21128 45404
rect 20947 45373 20959 45376
rect 20901 45367 20959 45373
rect 21100 45348 21128 45376
rect 22281 45373 22293 45407
rect 22327 45404 22339 45407
rect 22922 45404 22928 45416
rect 22327 45376 22928 45404
rect 22327 45373 22339 45376
rect 22281 45367 22339 45373
rect 22922 45364 22928 45376
rect 22980 45364 22986 45416
rect 12897 45339 12955 45345
rect 12897 45305 12909 45339
rect 12943 45336 12955 45339
rect 13906 45336 13912 45348
rect 12943 45308 13912 45336
rect 12943 45305 12955 45308
rect 12897 45299 12955 45305
rect 13906 45296 13912 45308
rect 13964 45296 13970 45348
rect 19153 45339 19211 45345
rect 19153 45305 19165 45339
rect 19199 45336 19211 45339
rect 19334 45336 19340 45348
rect 19199 45308 19340 45336
rect 19199 45305 19211 45308
rect 19153 45299 19211 45305
rect 19334 45296 19340 45308
rect 19392 45296 19398 45348
rect 21082 45296 21088 45348
rect 21140 45296 21146 45348
rect 29917 45339 29975 45345
rect 29917 45336 29929 45339
rect 22066 45308 29929 45336
rect 15470 45228 15476 45280
rect 15528 45268 15534 45280
rect 22066 45268 22094 45308
rect 29917 45305 29929 45308
rect 29963 45305 29975 45339
rect 29917 45299 29975 45305
rect 22922 45268 22928 45280
rect 15528 45240 22094 45268
rect 22883 45240 22928 45268
rect 15528 45228 15534 45240
rect 22922 45228 22928 45240
rect 22980 45228 22986 45280
rect 1104 45178 38824 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 38824 45178
rect 1104 45104 38824 45126
rect 21358 45064 21364 45076
rect 21319 45036 21364 45064
rect 21358 45024 21364 45036
rect 21416 45024 21422 45076
rect 17494 44956 17500 45008
rect 17552 44996 17558 45008
rect 25038 44996 25044 45008
rect 17552 44968 25044 44996
rect 17552 44956 17558 44968
rect 25038 44956 25044 44968
rect 25096 44956 25102 45008
rect 17865 44931 17923 44937
rect 17865 44897 17877 44931
rect 17911 44928 17923 44931
rect 18690 44928 18696 44940
rect 17911 44900 18696 44928
rect 17911 44897 17923 44900
rect 17865 44891 17923 44897
rect 18690 44888 18696 44900
rect 18748 44888 18754 44940
rect 19613 44931 19671 44937
rect 19613 44897 19625 44931
rect 19659 44928 19671 44931
rect 19978 44928 19984 44940
rect 19659 44900 19984 44928
rect 19659 44897 19671 44900
rect 19613 44891 19671 44897
rect 19978 44888 19984 44900
rect 20036 44888 20042 44940
rect 22462 44888 22468 44940
rect 22520 44928 22526 44940
rect 23293 44931 23351 44937
rect 23293 44928 23305 44931
rect 22520 44900 23305 44928
rect 22520 44888 22526 44900
rect 23293 44897 23305 44900
rect 23339 44897 23351 44931
rect 23293 44891 23351 44897
rect 18138 44860 18144 44872
rect 18099 44832 18144 44860
rect 18138 44820 18144 44832
rect 18196 44820 18202 44872
rect 19242 44820 19248 44872
rect 19300 44860 19306 44872
rect 19337 44863 19395 44869
rect 19337 44860 19349 44863
rect 19300 44832 19349 44860
rect 19300 44820 19306 44832
rect 19337 44829 19349 44832
rect 19383 44829 19395 44863
rect 23014 44860 23020 44872
rect 22975 44832 23020 44860
rect 19337 44823 19395 44829
rect 23014 44820 23020 44832
rect 23072 44820 23078 44872
rect 21269 44795 21327 44801
rect 21269 44761 21281 44795
rect 21315 44792 21327 44795
rect 21726 44792 21732 44804
rect 21315 44764 21732 44792
rect 21315 44761 21327 44764
rect 21269 44755 21327 44761
rect 21726 44752 21732 44764
rect 21784 44752 21790 44804
rect 1104 44634 38824 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 38824 44634
rect 1104 44560 38824 44582
rect 16117 44523 16175 44529
rect 16117 44489 16129 44523
rect 16163 44520 16175 44523
rect 16850 44520 16856 44532
rect 16163 44492 16856 44520
rect 16163 44489 16175 44492
rect 16117 44483 16175 44489
rect 16850 44480 16856 44492
rect 16908 44520 16914 44532
rect 17310 44520 17316 44532
rect 16908 44492 17316 44520
rect 16908 44480 16914 44492
rect 17310 44480 17316 44492
rect 17368 44480 17374 44532
rect 18322 44520 18328 44532
rect 18283 44492 18328 44520
rect 18322 44480 18328 44492
rect 18380 44480 18386 44532
rect 23845 44523 23903 44529
rect 23845 44489 23857 44523
rect 23891 44520 23903 44523
rect 24394 44520 24400 44532
rect 23891 44492 24400 44520
rect 23891 44489 23903 44492
rect 23845 44483 23903 44489
rect 24394 44480 24400 44492
rect 24452 44480 24458 44532
rect 13164 44387 13222 44393
rect 13164 44353 13176 44387
rect 13210 44384 13222 44387
rect 14550 44384 14556 44396
rect 13210 44356 14556 44384
rect 13210 44353 13222 44356
rect 13164 44347 13222 44353
rect 14550 44344 14556 44356
rect 14608 44344 14614 44396
rect 14826 44344 14832 44396
rect 14884 44384 14890 44396
rect 14993 44387 15051 44393
rect 14993 44384 15005 44387
rect 14884 44356 15005 44384
rect 14884 44344 14890 44356
rect 14993 44353 15005 44356
rect 15039 44353 15051 44387
rect 14993 44347 15051 44353
rect 18046 44344 18052 44396
rect 18104 44384 18110 44396
rect 20070 44393 20076 44396
rect 18141 44387 18199 44393
rect 18141 44384 18153 44387
rect 18104 44356 18153 44384
rect 18104 44344 18110 44356
rect 18141 44353 18153 44356
rect 18187 44353 18199 44387
rect 18141 44347 18199 44353
rect 20064 44347 20076 44393
rect 20128 44384 20134 44396
rect 20128 44356 20164 44384
rect 20070 44344 20076 44347
rect 20128 44344 20134 44356
rect 20990 44344 20996 44396
rect 21048 44384 21054 44396
rect 22833 44387 22891 44393
rect 22833 44384 22845 44387
rect 21048 44356 22845 44384
rect 21048 44344 21054 44356
rect 22833 44353 22845 44356
rect 22879 44353 22891 44387
rect 24026 44384 24032 44396
rect 23987 44356 24032 44384
rect 22833 44347 22891 44353
rect 24026 44344 24032 44356
rect 24084 44344 24090 44396
rect 12894 44316 12900 44328
rect 12855 44288 12900 44316
rect 12894 44276 12900 44288
rect 12952 44276 12958 44328
rect 14642 44276 14648 44328
rect 14700 44316 14706 44328
rect 14737 44319 14795 44325
rect 14737 44316 14749 44319
rect 14700 44288 14749 44316
rect 14700 44276 14706 44288
rect 14737 44285 14749 44288
rect 14783 44285 14795 44319
rect 14737 44279 14795 44285
rect 17957 44319 18015 44325
rect 17957 44285 17969 44319
rect 18003 44316 18015 44319
rect 19794 44316 19800 44328
rect 18003 44288 18184 44316
rect 19755 44288 19800 44316
rect 18003 44285 18015 44288
rect 17957 44279 18015 44285
rect 18156 44260 18184 44288
rect 19794 44276 19800 44288
rect 19852 44276 19858 44328
rect 22557 44319 22615 44325
rect 22557 44285 22569 44319
rect 22603 44316 22615 44319
rect 23474 44316 23480 44328
rect 22603 44288 23480 44316
rect 22603 44285 22615 44288
rect 22557 44279 22615 44285
rect 23474 44276 23480 44288
rect 23532 44276 23538 44328
rect 18138 44208 18144 44260
rect 18196 44208 18202 44260
rect 14277 44183 14335 44189
rect 14277 44149 14289 44183
rect 14323 44180 14335 44183
rect 14458 44180 14464 44192
rect 14323 44152 14464 44180
rect 14323 44149 14335 44152
rect 14277 44143 14335 44149
rect 14458 44140 14464 44152
rect 14516 44140 14522 44192
rect 21082 44140 21088 44192
rect 21140 44180 21146 44192
rect 21177 44183 21235 44189
rect 21177 44180 21189 44183
rect 21140 44152 21189 44180
rect 21140 44140 21146 44152
rect 21177 44149 21189 44152
rect 21223 44149 21235 44183
rect 21177 44143 21235 44149
rect 1104 44090 38824 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 38824 44090
rect 1104 44016 38824 44038
rect 19978 43936 19984 43988
rect 20036 43976 20042 43988
rect 20622 43976 20628 43988
rect 20036 43948 20628 43976
rect 20036 43936 20042 43948
rect 20622 43936 20628 43948
rect 20680 43936 20686 43988
rect 22646 43976 22652 43988
rect 20732 43948 22652 43976
rect 20254 43868 20260 43920
rect 20312 43908 20318 43920
rect 20732 43908 20760 43948
rect 22646 43936 22652 43948
rect 22704 43936 22710 43988
rect 23293 43979 23351 43985
rect 23293 43945 23305 43979
rect 23339 43976 23351 43979
rect 24026 43976 24032 43988
rect 23339 43948 24032 43976
rect 23339 43945 23351 43948
rect 23293 43939 23351 43945
rect 24026 43936 24032 43948
rect 24084 43936 24090 43988
rect 20312 43880 20760 43908
rect 20312 43868 20318 43880
rect 17773 43843 17831 43849
rect 17773 43809 17785 43843
rect 17819 43840 17831 43843
rect 18046 43840 18052 43852
rect 17819 43812 18052 43840
rect 17819 43809 17831 43812
rect 17773 43803 17831 43809
rect 18046 43800 18052 43812
rect 18104 43800 18110 43852
rect 14277 43775 14335 43781
rect 14277 43741 14289 43775
rect 14323 43772 14335 43775
rect 14458 43772 14464 43784
rect 14323 43744 14464 43772
rect 14323 43741 14335 43744
rect 14277 43735 14335 43741
rect 14458 43732 14464 43744
rect 14516 43732 14522 43784
rect 14642 43732 14648 43784
rect 14700 43772 14706 43784
rect 15657 43775 15715 43781
rect 15657 43772 15669 43775
rect 14700 43744 15669 43772
rect 14700 43732 14706 43744
rect 15657 43741 15669 43744
rect 15703 43772 15715 43775
rect 16666 43772 16672 43784
rect 15703 43744 16672 43772
rect 15703 43741 15715 43744
rect 15657 43735 15715 43741
rect 16666 43732 16672 43744
rect 16724 43732 16730 43784
rect 17494 43772 17500 43784
rect 17455 43744 17500 43772
rect 17494 43732 17500 43744
rect 17552 43732 17558 43784
rect 19245 43775 19303 43781
rect 19245 43741 19257 43775
rect 19291 43772 19303 43775
rect 19794 43772 19800 43784
rect 19291 43744 19800 43772
rect 19291 43741 19303 43744
rect 19245 43735 19303 43741
rect 19794 43732 19800 43744
rect 19852 43772 19858 43784
rect 20901 43775 20959 43781
rect 20901 43772 20913 43775
rect 19852 43744 20913 43772
rect 19852 43732 19858 43744
rect 20901 43741 20913 43744
rect 20947 43772 20959 43775
rect 22002 43772 22008 43784
rect 20947 43744 22008 43772
rect 20947 43741 20959 43744
rect 20901 43735 20959 43741
rect 22002 43732 22008 43744
rect 22060 43732 22066 43784
rect 22925 43775 22983 43781
rect 22925 43772 22937 43775
rect 22296 43744 22937 43772
rect 14093 43707 14151 43713
rect 14093 43673 14105 43707
rect 14139 43704 14151 43707
rect 14139 43676 15148 43704
rect 14139 43673 14151 43676
rect 14093 43667 14151 43673
rect 14461 43639 14519 43645
rect 14461 43605 14473 43639
rect 14507 43636 14519 43639
rect 15010 43636 15016 43648
rect 14507 43608 15016 43636
rect 14507 43605 14519 43608
rect 14461 43599 14519 43605
rect 15010 43596 15016 43608
rect 15068 43596 15074 43648
rect 15120 43636 15148 43676
rect 15286 43664 15292 43716
rect 15344 43704 15350 43716
rect 15902 43707 15960 43713
rect 15902 43704 15914 43707
rect 15344 43676 15914 43704
rect 15344 43664 15350 43676
rect 15902 43673 15914 43676
rect 15948 43673 15960 43707
rect 15902 43667 15960 43673
rect 19334 43664 19340 43716
rect 19392 43704 19398 43716
rect 19490 43707 19548 43713
rect 19490 43704 19502 43707
rect 19392 43676 19502 43704
rect 19392 43664 19398 43676
rect 19490 43673 19502 43676
rect 19536 43673 19548 43707
rect 19490 43667 19548 43673
rect 20714 43664 20720 43716
rect 20772 43704 20778 43716
rect 21146 43707 21204 43713
rect 21146 43704 21158 43707
rect 20772 43676 21158 43704
rect 20772 43664 20778 43676
rect 21146 43673 21158 43676
rect 21192 43673 21204 43707
rect 21146 43667 21204 43673
rect 15378 43636 15384 43648
rect 15120 43608 15384 43636
rect 15378 43596 15384 43608
rect 15436 43596 15442 43648
rect 17037 43639 17095 43645
rect 17037 43605 17049 43639
rect 17083 43636 17095 43639
rect 17218 43636 17224 43648
rect 17083 43608 17224 43636
rect 17083 43605 17095 43608
rect 17037 43599 17095 43605
rect 17218 43596 17224 43608
rect 17276 43596 17282 43648
rect 22094 43596 22100 43648
rect 22152 43636 22158 43648
rect 22296 43645 22324 43744
rect 22925 43741 22937 43744
rect 22971 43741 22983 43775
rect 22925 43735 22983 43741
rect 23109 43775 23167 43781
rect 23109 43741 23121 43775
rect 23155 43772 23167 43775
rect 23290 43772 23296 43784
rect 23155 43744 23296 43772
rect 23155 43741 23167 43744
rect 23109 43735 23167 43741
rect 22646 43704 22652 43716
rect 22559 43676 22652 43704
rect 22646 43664 22652 43676
rect 22704 43704 22710 43716
rect 23124 43704 23152 43735
rect 23290 43732 23296 43744
rect 23348 43732 23354 43784
rect 22704 43676 23152 43704
rect 22704 43664 22710 43676
rect 22281 43639 22339 43645
rect 22281 43636 22293 43639
rect 22152 43608 22293 43636
rect 22152 43596 22158 43608
rect 22281 43605 22293 43608
rect 22327 43605 22339 43639
rect 22281 43599 22339 43605
rect 1104 43546 38824 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 38824 43546
rect 1104 43472 38824 43494
rect 14090 43432 14096 43444
rect 14051 43404 14096 43432
rect 14090 43392 14096 43404
rect 14148 43392 14154 43444
rect 14550 43432 14556 43444
rect 14511 43404 14556 43432
rect 14550 43392 14556 43404
rect 14608 43392 14614 43444
rect 23934 43432 23940 43444
rect 23895 43404 23940 43432
rect 23934 43392 23940 43404
rect 23992 43392 23998 43444
rect 24578 43432 24584 43444
rect 24539 43404 24584 43432
rect 24578 43392 24584 43404
rect 24636 43392 24642 43444
rect 14642 43364 14648 43376
rect 12728 43336 14648 43364
rect 12728 43305 12756 43336
rect 14642 43324 14648 43336
rect 14700 43324 14706 43376
rect 20073 43367 20131 43373
rect 20073 43333 20085 43367
rect 20119 43364 20131 43367
rect 21082 43364 21088 43376
rect 20119 43336 21088 43364
rect 20119 43333 20131 43336
rect 20073 43327 20131 43333
rect 21082 43324 21088 43336
rect 21140 43324 21146 43376
rect 12713 43299 12771 43305
rect 12713 43265 12725 43299
rect 12759 43265 12771 43299
rect 12713 43259 12771 43265
rect 12980 43299 13038 43305
rect 12980 43265 12992 43299
rect 13026 43296 13038 43299
rect 14090 43296 14096 43308
rect 13026 43268 14096 43296
rect 13026 43265 13038 43268
rect 12980 43259 13038 43265
rect 14090 43256 14096 43268
rect 14148 43256 14154 43308
rect 14783 43299 14841 43305
rect 14783 43296 14795 43299
rect 14660 43268 14795 43296
rect 14660 43160 14688 43268
rect 14783 43265 14795 43268
rect 14829 43265 14841 43299
rect 14918 43296 14924 43308
rect 14879 43268 14924 43296
rect 14783 43259 14841 43265
rect 14918 43256 14924 43268
rect 14976 43256 14982 43308
rect 15010 43256 15016 43308
rect 15068 43296 15074 43308
rect 15194 43296 15200 43308
rect 15068 43268 15113 43296
rect 15155 43268 15200 43296
rect 15068 43256 15074 43268
rect 15194 43256 15200 43268
rect 15252 43256 15258 43308
rect 15378 43256 15384 43308
rect 15436 43296 15442 43308
rect 15749 43299 15807 43305
rect 15749 43296 15761 43299
rect 15436 43268 15761 43296
rect 15436 43256 15442 43268
rect 15749 43265 15761 43268
rect 15795 43265 15807 43299
rect 15749 43259 15807 43265
rect 15933 43299 15991 43305
rect 15933 43265 15945 43299
rect 15979 43296 15991 43299
rect 16666 43296 16672 43308
rect 15979 43268 16528 43296
rect 16627 43268 16672 43296
rect 15979 43265 15991 43268
rect 15933 43259 15991 43265
rect 15930 43160 15936 43172
rect 14660 43132 15936 43160
rect 15930 43120 15936 43132
rect 15988 43120 15994 43172
rect 16022 43052 16028 43104
rect 16080 43092 16086 43104
rect 16117 43095 16175 43101
rect 16117 43092 16129 43095
rect 16080 43064 16129 43092
rect 16080 43052 16086 43064
rect 16117 43061 16129 43064
rect 16163 43061 16175 43095
rect 16500 43092 16528 43268
rect 16666 43256 16672 43268
rect 16724 43256 16730 43308
rect 16758 43256 16764 43308
rect 16816 43296 16822 43308
rect 16925 43299 16983 43305
rect 16925 43296 16937 43299
rect 16816 43268 16937 43296
rect 16816 43256 16822 43268
rect 16925 43265 16937 43268
rect 16971 43265 16983 43299
rect 19886 43296 19892 43308
rect 19847 43268 19892 43296
rect 16925 43259 16983 43265
rect 19886 43256 19892 43268
rect 19944 43256 19950 43308
rect 24118 43296 24124 43308
rect 24079 43268 24124 43296
rect 24118 43256 24124 43268
rect 24176 43256 24182 43308
rect 24762 43296 24768 43308
rect 24723 43268 24768 43296
rect 24762 43256 24768 43268
rect 24820 43256 24826 43308
rect 18049 43095 18107 43101
rect 18049 43092 18061 43095
rect 16500 43064 18061 43092
rect 16117 43055 16175 43061
rect 18049 43061 18061 43064
rect 18095 43092 18107 43095
rect 18138 43092 18144 43104
rect 18095 43064 18144 43092
rect 18095 43061 18107 43064
rect 18049 43055 18107 43061
rect 18138 43052 18144 43064
rect 18196 43052 18202 43104
rect 20257 43095 20315 43101
rect 20257 43061 20269 43095
rect 20303 43092 20315 43095
rect 20622 43092 20628 43104
rect 20303 43064 20628 43092
rect 20303 43061 20315 43064
rect 20257 43055 20315 43061
rect 20622 43052 20628 43064
rect 20680 43052 20686 43104
rect 1104 43002 38824 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 38824 43002
rect 1104 42928 38824 42950
rect 15565 42891 15623 42897
rect 15565 42857 15577 42891
rect 15611 42888 15623 42891
rect 16758 42888 16764 42900
rect 15611 42860 16764 42888
rect 15611 42857 15623 42860
rect 15565 42851 15623 42857
rect 16758 42848 16764 42860
rect 16816 42848 16822 42900
rect 24762 42888 24768 42900
rect 24723 42860 24768 42888
rect 24762 42848 24768 42860
rect 24820 42848 24826 42900
rect 20533 42823 20591 42829
rect 20533 42789 20545 42823
rect 20579 42820 20591 42823
rect 20714 42820 20720 42832
rect 20579 42792 20720 42820
rect 20579 42789 20591 42792
rect 20533 42783 20591 42789
rect 20714 42780 20720 42792
rect 20772 42780 20778 42832
rect 20898 42780 20904 42832
rect 20956 42780 20962 42832
rect 14090 42752 14096 42764
rect 14051 42724 14096 42752
rect 14090 42712 14096 42724
rect 14148 42712 14154 42764
rect 14182 42712 14188 42764
rect 14240 42752 14246 42764
rect 14918 42752 14924 42764
rect 14240 42724 14924 42752
rect 14240 42712 14246 42724
rect 13357 42687 13415 42693
rect 13357 42653 13369 42687
rect 13403 42684 13415 42687
rect 13998 42684 14004 42696
rect 13403 42656 14004 42684
rect 13403 42653 13415 42656
rect 13357 42647 13415 42653
rect 13998 42644 14004 42656
rect 14056 42644 14062 42696
rect 14366 42684 14372 42696
rect 14327 42656 14372 42684
rect 14366 42644 14372 42656
rect 14424 42644 14430 42696
rect 14476 42693 14504 42724
rect 14918 42712 14924 42724
rect 14976 42752 14982 42764
rect 14976 42724 15976 42752
rect 14976 42712 14982 42724
rect 14461 42687 14519 42693
rect 14461 42653 14473 42687
rect 14507 42653 14519 42687
rect 14461 42647 14519 42653
rect 14553 42687 14611 42693
rect 14553 42653 14565 42687
rect 14599 42653 14611 42687
rect 14734 42684 14740 42696
rect 14695 42656 14740 42684
rect 14553 42647 14611 42653
rect 13173 42619 13231 42625
rect 13173 42585 13185 42619
rect 13219 42616 13231 42619
rect 13262 42616 13268 42628
rect 13219 42588 13268 42616
rect 13219 42585 13231 42588
rect 13173 42579 13231 42585
rect 13262 42576 13268 42588
rect 13320 42576 13326 42628
rect 13541 42619 13599 42625
rect 13541 42585 13553 42619
rect 13587 42616 13599 42619
rect 14568 42616 14596 42647
rect 14734 42644 14740 42656
rect 14792 42684 14798 42696
rect 15194 42684 15200 42696
rect 14792 42656 15200 42684
rect 14792 42644 14798 42656
rect 15194 42644 15200 42656
rect 15252 42644 15258 42696
rect 15948 42693 15976 42724
rect 15841 42687 15899 42693
rect 15841 42653 15853 42687
rect 15887 42653 15899 42687
rect 15841 42647 15899 42653
rect 15933 42687 15991 42693
rect 15933 42653 15945 42687
rect 15979 42653 15991 42687
rect 15933 42647 15991 42653
rect 13587 42588 14596 42616
rect 15856 42616 15884 42647
rect 16022 42644 16028 42696
rect 16080 42684 16086 42696
rect 16080 42656 16125 42684
rect 16080 42644 16086 42656
rect 16206 42644 16212 42696
rect 16264 42684 16270 42696
rect 19521 42687 19579 42693
rect 16264 42656 16309 42684
rect 16264 42644 16270 42656
rect 19521 42653 19533 42687
rect 19567 42684 19579 42687
rect 19978 42684 19984 42696
rect 19567 42656 19984 42684
rect 19567 42653 19579 42656
rect 19521 42647 19579 42653
rect 19978 42644 19984 42656
rect 20036 42684 20042 42696
rect 20254 42684 20260 42696
rect 20036 42656 20260 42684
rect 20036 42644 20042 42656
rect 20254 42644 20260 42656
rect 20312 42644 20318 42696
rect 20913 42693 20941 42780
rect 22005 42755 22063 42761
rect 22005 42752 22017 42755
rect 21021 42724 22017 42752
rect 21021 42693 21049 42724
rect 22005 42721 22017 42724
rect 22051 42721 22063 42755
rect 22005 42715 22063 42721
rect 23382 42712 23388 42764
rect 23440 42752 23446 42764
rect 25041 42755 25099 42761
rect 25041 42752 25053 42755
rect 23440 42724 25053 42752
rect 23440 42712 23446 42724
rect 20809 42687 20867 42693
rect 20809 42653 20821 42687
rect 20855 42653 20867 42687
rect 20809 42647 20867 42653
rect 20898 42687 20956 42693
rect 20898 42653 20910 42687
rect 20944 42653 20956 42687
rect 20898 42647 20956 42653
rect 21014 42687 21072 42693
rect 21014 42653 21026 42687
rect 21060 42653 21072 42687
rect 21174 42684 21180 42696
rect 21135 42656 21180 42684
rect 21014 42647 21072 42653
rect 17402 42616 17408 42628
rect 15856 42588 17408 42616
rect 13587 42585 13599 42588
rect 13541 42579 13599 42585
rect 17402 42576 17408 42588
rect 17460 42576 17466 42628
rect 19337 42619 19395 42625
rect 19337 42585 19349 42619
rect 19383 42616 19395 42619
rect 19886 42616 19892 42628
rect 19383 42588 19892 42616
rect 19383 42585 19395 42588
rect 19337 42579 19395 42585
rect 19886 42576 19892 42588
rect 19944 42616 19950 42628
rect 19944 42588 20116 42616
rect 19944 42576 19950 42588
rect 13998 42508 14004 42560
rect 14056 42548 14062 42560
rect 14918 42548 14924 42560
rect 14056 42520 14924 42548
rect 14056 42508 14062 42520
rect 14918 42508 14924 42520
rect 14976 42508 14982 42560
rect 19426 42508 19432 42560
rect 19484 42548 19490 42560
rect 19705 42551 19763 42557
rect 19705 42548 19717 42551
rect 19484 42520 19717 42548
rect 19484 42508 19490 42520
rect 19705 42517 19717 42520
rect 19751 42517 19763 42551
rect 20088 42548 20116 42588
rect 20714 42576 20720 42628
rect 20772 42616 20778 42628
rect 20824 42616 20852 42647
rect 21174 42644 21180 42656
rect 21232 42644 21238 42696
rect 24596 42693 24624 42724
rect 25041 42721 25053 42724
rect 25087 42752 25099 42755
rect 27706 42752 27712 42764
rect 25087 42724 27712 42752
rect 25087 42721 25099 42724
rect 25041 42715 25099 42721
rect 27706 42712 27712 42724
rect 27764 42712 27770 42764
rect 24397 42687 24455 42693
rect 24397 42653 24409 42687
rect 24443 42653 24455 42687
rect 24397 42647 24455 42653
rect 24581 42687 24639 42693
rect 24581 42653 24593 42687
rect 24627 42653 24639 42687
rect 24581 42647 24639 42653
rect 20772 42588 20852 42616
rect 21637 42619 21695 42625
rect 20772 42576 20778 42588
rect 21637 42585 21649 42619
rect 21683 42585 21695 42619
rect 21637 42579 21695 42585
rect 21821 42619 21879 42625
rect 21821 42585 21833 42619
rect 21867 42616 21879 42619
rect 22094 42616 22100 42628
rect 21867 42588 22100 42616
rect 21867 42585 21879 42588
rect 21821 42579 21879 42585
rect 20438 42548 20444 42560
rect 20088 42520 20444 42548
rect 19705 42511 19763 42517
rect 20438 42508 20444 42520
rect 20496 42548 20502 42560
rect 21652 42548 21680 42579
rect 22094 42576 22100 42588
rect 22152 42576 22158 42628
rect 22465 42619 22523 42625
rect 22465 42585 22477 42619
rect 22511 42585 22523 42619
rect 22646 42616 22652 42628
rect 22607 42588 22652 42616
rect 22465 42579 22523 42585
rect 22480 42548 22508 42579
rect 22646 42576 22652 42588
rect 22704 42616 22710 42628
rect 24412 42616 24440 42647
rect 22704 42588 24440 42616
rect 22704 42576 22710 42588
rect 22830 42548 22836 42560
rect 20496 42520 22508 42548
rect 22791 42520 22836 42548
rect 20496 42508 20502 42520
rect 22830 42508 22836 42520
rect 22888 42508 22894 42560
rect 1104 42458 38824 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 38824 42458
rect 1104 42384 38824 42406
rect 14185 42347 14243 42353
rect 14185 42313 14197 42347
rect 14231 42344 14243 42347
rect 14826 42344 14832 42356
rect 14231 42316 14832 42344
rect 14231 42313 14243 42316
rect 14185 42307 14243 42313
rect 14826 42304 14832 42316
rect 14884 42304 14890 42356
rect 15286 42344 15292 42356
rect 15247 42316 15292 42344
rect 15286 42304 15292 42316
rect 15344 42304 15350 42356
rect 17494 42344 17500 42356
rect 17455 42316 17500 42344
rect 17494 42304 17500 42316
rect 17552 42304 17558 42356
rect 19061 42347 19119 42353
rect 19061 42313 19073 42347
rect 19107 42344 19119 42347
rect 19334 42344 19340 42356
rect 19107 42316 19340 42344
rect 19107 42313 19119 42316
rect 19061 42307 19119 42313
rect 19334 42304 19340 42316
rect 19392 42304 19398 42356
rect 20070 42304 20076 42356
rect 20128 42344 20134 42356
rect 20165 42347 20223 42353
rect 20165 42344 20177 42347
rect 20128 42316 20177 42344
rect 20128 42304 20134 42316
rect 20165 42313 20177 42316
rect 20211 42313 20223 42347
rect 20165 42307 20223 42313
rect 24118 42304 24124 42356
rect 24176 42344 24182 42356
rect 24213 42347 24271 42353
rect 24213 42344 24225 42347
rect 24176 42316 24225 42344
rect 24176 42304 24182 42316
rect 24213 42313 24225 42316
rect 24259 42313 24271 42347
rect 24213 42307 24271 42313
rect 16298 42276 16304 42288
rect 14660 42248 16304 42276
rect 14274 42168 14280 42220
rect 14332 42208 14338 42220
rect 14660 42217 14688 42248
rect 16298 42236 16304 42248
rect 16356 42236 16362 42288
rect 20898 42276 20904 42288
rect 19444 42248 20904 42276
rect 14415 42211 14473 42217
rect 14415 42208 14427 42211
rect 14332 42180 14427 42208
rect 14332 42168 14338 42180
rect 14415 42177 14427 42180
rect 14461 42177 14473 42211
rect 14415 42171 14473 42177
rect 14566 42211 14624 42217
rect 14566 42177 14578 42211
rect 14612 42177 14624 42211
rect 14660 42211 14724 42217
rect 14660 42180 14678 42211
rect 14566 42171 14624 42177
rect 14666 42177 14678 42180
rect 14712 42177 14724 42211
rect 14826 42208 14832 42220
rect 14787 42180 14832 42208
rect 14666 42171 14724 42177
rect 14182 42100 14188 42152
rect 14240 42140 14246 42152
rect 14568 42140 14596 42171
rect 14826 42168 14832 42180
rect 14884 42168 14890 42220
rect 15562 42217 15568 42220
rect 15519 42211 15568 42217
rect 15519 42177 15531 42211
rect 15565 42177 15568 42211
rect 15519 42171 15568 42177
rect 15562 42168 15568 42171
rect 15620 42168 15626 42220
rect 15654 42211 15712 42217
rect 15654 42177 15666 42211
rect 15700 42177 15712 42211
rect 15654 42171 15712 42177
rect 15749 42211 15807 42217
rect 15749 42177 15761 42211
rect 15795 42208 15807 42211
rect 15838 42208 15844 42220
rect 15795 42180 15844 42208
rect 15795 42177 15807 42180
rect 15749 42171 15807 42177
rect 14240 42112 14596 42140
rect 14240 42100 14246 42112
rect 14568 42072 14596 42112
rect 15672 42072 15700 42171
rect 15838 42168 15844 42180
rect 15896 42168 15902 42220
rect 15933 42211 15991 42217
rect 15933 42177 15945 42211
rect 15979 42208 15991 42211
rect 16114 42208 16120 42220
rect 15979 42180 16120 42208
rect 15979 42177 15991 42180
rect 15933 42171 15991 42177
rect 14568 42044 15700 42072
rect 14366 41964 14372 42016
rect 14424 42004 14430 42016
rect 14734 42004 14740 42016
rect 14424 41976 14740 42004
rect 14424 41964 14430 41976
rect 14734 41964 14740 41976
rect 14792 41964 14798 42016
rect 14826 41964 14832 42016
rect 14884 42004 14890 42016
rect 15948 42004 15976 42171
rect 16114 42168 16120 42180
rect 16172 42168 16178 42220
rect 18046 42168 18052 42220
rect 18104 42208 18110 42220
rect 19444 42217 19472 42248
rect 18141 42211 18199 42217
rect 18141 42208 18153 42211
rect 18104 42180 18153 42208
rect 18104 42168 18110 42180
rect 18141 42177 18153 42180
rect 18187 42177 18199 42211
rect 18141 42171 18199 42177
rect 19291 42211 19349 42217
rect 19291 42177 19303 42211
rect 19337 42177 19349 42211
rect 19291 42171 19349 42177
rect 19429 42211 19487 42217
rect 19429 42177 19441 42211
rect 19475 42177 19487 42211
rect 19429 42171 19487 42177
rect 16206 42100 16212 42152
rect 16264 42140 16270 42152
rect 17037 42143 17095 42149
rect 17037 42140 17049 42143
rect 16264 42112 17049 42140
rect 16264 42100 16270 42112
rect 17037 42109 17049 42112
rect 17083 42109 17095 42143
rect 17037 42103 17095 42109
rect 17310 42072 17316 42084
rect 17271 42044 17316 42072
rect 17310 42032 17316 42044
rect 17368 42032 17374 42084
rect 19306 42072 19334 42171
rect 19518 42168 19524 42220
rect 19576 42208 19582 42220
rect 19705 42211 19763 42217
rect 19576 42180 19621 42208
rect 19576 42168 19582 42180
rect 19705 42177 19717 42211
rect 19751 42177 19763 42211
rect 19705 42171 19763 42177
rect 19720 42140 19748 42171
rect 20346 42168 20352 42220
rect 20404 42208 20410 42220
rect 20548 42217 20576 42248
rect 20898 42236 20904 42248
rect 20956 42236 20962 42288
rect 20441 42211 20499 42217
rect 20441 42208 20453 42211
rect 20404 42180 20453 42208
rect 20404 42168 20410 42180
rect 20441 42177 20453 42180
rect 20487 42177 20499 42211
rect 20441 42171 20499 42177
rect 20533 42211 20591 42217
rect 20533 42177 20545 42211
rect 20579 42177 20591 42211
rect 20533 42171 20591 42177
rect 20622 42168 20628 42220
rect 20680 42208 20686 42220
rect 20680 42180 20725 42208
rect 20680 42168 20686 42180
rect 20806 42168 20812 42220
rect 20864 42208 20870 42220
rect 21174 42208 21180 42220
rect 20864 42180 21180 42208
rect 20864 42168 20870 42180
rect 21174 42168 21180 42180
rect 21232 42168 21238 42220
rect 22002 42208 22008 42220
rect 21963 42180 22008 42208
rect 22002 42168 22008 42180
rect 22060 42168 22066 42220
rect 22261 42211 22319 42217
rect 22261 42208 22273 42211
rect 22112 42180 22273 42208
rect 20824 42140 20852 42168
rect 19720 42112 20852 42140
rect 21450 42100 21456 42152
rect 21508 42140 21514 42152
rect 22112 42140 22140 42180
rect 22261 42177 22273 42180
rect 22307 42177 22319 42211
rect 24026 42208 24032 42220
rect 23987 42180 24032 42208
rect 22261 42171 22319 42177
rect 24026 42168 24032 42180
rect 24084 42208 24090 42220
rect 27522 42208 27528 42220
rect 24084 42180 27528 42208
rect 24084 42168 24090 42180
rect 27522 42168 27528 42180
rect 27580 42168 27586 42220
rect 23842 42140 23848 42152
rect 21508 42112 22140 42140
rect 23803 42112 23848 42140
rect 21508 42100 21514 42112
rect 23842 42100 23848 42112
rect 23900 42100 23906 42152
rect 19978 42072 19984 42084
rect 19306 42044 19984 42072
rect 19978 42032 19984 42044
rect 20036 42032 20042 42084
rect 17954 42004 17960 42016
rect 14884 41976 15976 42004
rect 17915 41976 17960 42004
rect 14884 41964 14890 41976
rect 17954 41964 17960 41976
rect 18012 41964 18018 42016
rect 20254 41964 20260 42016
rect 20312 42004 20318 42016
rect 20438 42004 20444 42016
rect 20312 41976 20444 42004
rect 20312 41964 20318 41976
rect 20438 41964 20444 41976
rect 20496 41964 20502 42016
rect 22646 41964 22652 42016
rect 22704 42004 22710 42016
rect 23385 42007 23443 42013
rect 23385 42004 23397 42007
rect 22704 41976 23397 42004
rect 22704 41964 22710 41976
rect 23385 41973 23397 41976
rect 23431 41973 23443 42007
rect 23385 41967 23443 41973
rect 1104 41914 38824 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 38824 41914
rect 1104 41840 38824 41862
rect 11514 41760 11520 41812
rect 11572 41800 11578 41812
rect 11572 41772 12434 41800
rect 11572 41760 11578 41772
rect 12406 41732 12434 41772
rect 16666 41760 16672 41812
rect 16724 41800 16730 41812
rect 17129 41803 17187 41809
rect 17129 41800 17141 41803
rect 16724 41772 17141 41800
rect 16724 41760 16730 41772
rect 17129 41769 17141 41772
rect 17175 41800 17187 41803
rect 17678 41800 17684 41812
rect 17175 41772 17684 41800
rect 17175 41769 17187 41772
rect 17129 41763 17187 41769
rect 17678 41760 17684 41772
rect 17736 41760 17742 41812
rect 22002 41760 22008 41812
rect 22060 41800 22066 41812
rect 22557 41803 22615 41809
rect 22557 41800 22569 41803
rect 22060 41772 22569 41800
rect 22060 41760 22066 41772
rect 22557 41769 22569 41772
rect 22603 41769 22615 41803
rect 27522 41800 27528 41812
rect 27483 41772 27528 41800
rect 22557 41763 22615 41769
rect 27522 41760 27528 41772
rect 27580 41760 27586 41812
rect 24026 41732 24032 41744
rect 12406 41704 24032 41732
rect 24026 41692 24032 41704
rect 24084 41692 24090 41744
rect 14182 41624 14188 41676
rect 14240 41664 14246 41676
rect 14369 41667 14427 41673
rect 14369 41664 14381 41667
rect 14240 41636 14381 41664
rect 14240 41624 14246 41636
rect 14369 41633 14381 41636
rect 14415 41633 14427 41667
rect 14369 41627 14427 41633
rect 15286 41624 15292 41676
rect 15344 41664 15350 41676
rect 15838 41664 15844 41676
rect 15344 41636 15844 41664
rect 15344 41624 15350 41636
rect 15838 41624 15844 41636
rect 15896 41624 15902 41676
rect 13541 41599 13599 41605
rect 13541 41565 13553 41599
rect 13587 41565 13599 41599
rect 13541 41559 13599 41565
rect 14093 41599 14151 41605
rect 14093 41565 14105 41599
rect 14139 41596 14151 41599
rect 19613 41599 19671 41605
rect 19613 41596 19625 41599
rect 14139 41568 19625 41596
rect 14139 41565 14151 41568
rect 14093 41559 14151 41565
rect 13262 41420 13268 41472
rect 13320 41460 13326 41472
rect 13357 41463 13415 41469
rect 13357 41460 13369 41463
rect 13320 41432 13369 41460
rect 13320 41420 13326 41432
rect 13357 41429 13369 41432
rect 13403 41429 13415 41463
rect 13357 41423 13415 41429
rect 13446 41420 13452 41472
rect 13504 41460 13510 41472
rect 13556 41460 13584 41559
rect 14568 41540 14596 41568
rect 19613 41565 19625 41568
rect 19659 41565 19671 41599
rect 19613 41559 19671 41565
rect 19889 41599 19947 41605
rect 19889 41565 19901 41599
rect 19935 41596 19947 41599
rect 20898 41596 20904 41608
rect 19935 41568 20904 41596
rect 19935 41565 19947 41568
rect 19889 41559 19947 41565
rect 20898 41556 20904 41568
rect 20956 41596 20962 41608
rect 21174 41596 21180 41608
rect 20956 41568 21180 41596
rect 20956 41556 20962 41568
rect 21174 41556 21180 41568
rect 21232 41556 21238 41608
rect 14550 41488 14556 41540
rect 14608 41488 14614 41540
rect 15194 41488 15200 41540
rect 15252 41528 15258 41540
rect 15841 41531 15899 41537
rect 15841 41528 15853 41531
rect 15252 41500 15853 41528
rect 15252 41488 15258 41500
rect 15841 41497 15853 41500
rect 15887 41497 15899 41531
rect 15841 41491 15899 41497
rect 21269 41531 21327 41537
rect 21269 41497 21281 41531
rect 21315 41528 21327 41531
rect 27246 41528 27252 41540
rect 21315 41500 27252 41528
rect 21315 41497 21327 41500
rect 21269 41491 21327 41497
rect 27246 41488 27252 41500
rect 27304 41488 27310 41540
rect 27433 41531 27491 41537
rect 27433 41497 27445 41531
rect 27479 41528 27491 41531
rect 27982 41528 27988 41540
rect 27479 41500 27988 41528
rect 27479 41497 27491 41500
rect 27433 41491 27491 41497
rect 27982 41488 27988 41500
rect 28040 41488 28046 41540
rect 19334 41460 19340 41472
rect 13504 41432 19340 41460
rect 13504 41420 13510 41432
rect 19334 41420 19340 41432
rect 19392 41420 19398 41472
rect 1104 41370 38824 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 38824 41370
rect 1104 41296 38824 41318
rect 13262 41216 13268 41268
rect 13320 41256 13326 41268
rect 15105 41259 15163 41265
rect 13320 41228 14780 41256
rect 13320 41216 13326 41228
rect 12713 41191 12771 41197
rect 12713 41157 12725 41191
rect 12759 41157 12771 41191
rect 12713 41151 12771 41157
rect 12929 41191 12987 41197
rect 12929 41157 12941 41191
rect 12975 41188 12987 41191
rect 13170 41188 13176 41200
rect 12975 41160 13176 41188
rect 12975 41157 12987 41160
rect 12929 41151 12987 41157
rect 12728 41120 12756 41151
rect 13170 41148 13176 41160
rect 13228 41148 13234 41200
rect 14752 41197 14780 41228
rect 15105 41225 15117 41259
rect 15151 41256 15163 41259
rect 15286 41256 15292 41268
rect 15151 41228 15292 41256
rect 15151 41225 15163 41228
rect 15105 41219 15163 41225
rect 15286 41216 15292 41228
rect 15344 41216 15350 41268
rect 15473 41259 15531 41265
rect 15473 41225 15485 41259
rect 15519 41256 15531 41259
rect 15562 41256 15568 41268
rect 15519 41228 15568 41256
rect 15519 41225 15531 41228
rect 15473 41219 15531 41225
rect 15562 41216 15568 41228
rect 15620 41216 15626 41268
rect 16850 41256 16856 41268
rect 15672 41228 16856 41256
rect 14737 41191 14795 41197
rect 14737 41157 14749 41191
rect 14783 41188 14795 41191
rect 15378 41188 15384 41200
rect 14783 41160 15384 41188
rect 14783 41157 14795 41160
rect 14737 41151 14795 41157
rect 15378 41148 15384 41160
rect 15436 41148 15442 41200
rect 15672 41188 15700 41228
rect 16850 41216 16856 41228
rect 16908 41216 16914 41268
rect 17221 41259 17279 41265
rect 17221 41225 17233 41259
rect 17267 41256 17279 41259
rect 18046 41256 18052 41268
rect 17267 41228 18052 41256
rect 17267 41225 17279 41228
rect 17221 41219 17279 41225
rect 18046 41216 18052 41228
rect 18104 41216 18110 41268
rect 18322 41216 18328 41268
rect 18380 41256 18386 41268
rect 34054 41256 34060 41268
rect 18380 41228 34060 41256
rect 18380 41216 18386 41228
rect 34054 41216 34060 41228
rect 34112 41216 34118 41268
rect 15488 41160 15700 41188
rect 15749 41191 15807 41197
rect 13262 41120 13268 41132
rect 12728 41092 13268 41120
rect 13004 41064 13032 41092
rect 13262 41080 13268 41092
rect 13320 41080 13326 41132
rect 14921 41123 14979 41129
rect 14921 41089 14933 41123
rect 14967 41089 14979 41123
rect 15488 41120 15516 41160
rect 15749 41157 15761 41191
rect 15795 41188 15807 41191
rect 15838 41188 15844 41200
rect 15795 41160 15844 41188
rect 15795 41157 15807 41160
rect 15749 41151 15807 41157
rect 15838 41148 15844 41160
rect 15896 41148 15902 41200
rect 15965 41191 16023 41197
rect 15965 41157 15977 41191
rect 16011 41188 16023 41191
rect 16206 41188 16212 41200
rect 16011 41160 16212 41188
rect 16011 41157 16023 41160
rect 15965 41151 16023 41157
rect 16206 41148 16212 41160
rect 16264 41148 16270 41200
rect 17034 41188 17040 41200
rect 16995 41160 17040 41188
rect 17034 41148 17040 41160
rect 17092 41148 17098 41200
rect 17954 41197 17960 41200
rect 17948 41151 17960 41197
rect 18012 41188 18018 41200
rect 18012 41160 18048 41188
rect 17954 41148 17960 41151
rect 18012 41148 18018 41160
rect 18230 41148 18236 41200
rect 18288 41188 18294 41200
rect 21634 41188 21640 41200
rect 18288 41160 21640 41188
rect 18288 41148 18294 41160
rect 21634 41148 21640 41160
rect 21692 41148 21698 41200
rect 21818 41148 21824 41200
rect 21876 41188 21882 41200
rect 22158 41191 22216 41197
rect 22158 41188 22170 41191
rect 21876 41160 22170 41188
rect 21876 41148 21882 41160
rect 22158 41157 22170 41160
rect 22204 41157 22216 41191
rect 22158 41151 22216 41157
rect 22278 41148 22284 41200
rect 22336 41188 22342 41200
rect 34790 41188 34796 41200
rect 22336 41160 34796 41188
rect 22336 41148 22342 41160
rect 34790 41148 34796 41160
rect 34848 41148 34854 41200
rect 17678 41120 17684 41132
rect 14921 41083 14979 41089
rect 15212 41092 15516 41120
rect 17639 41092 17684 41120
rect 12986 41012 12992 41064
rect 13044 41012 13050 41064
rect 13541 41055 13599 41061
rect 13541 41021 13553 41055
rect 13587 41052 13599 41055
rect 13722 41052 13728 41064
rect 13587 41024 13728 41052
rect 13587 41021 13599 41024
rect 13541 41015 13599 41021
rect 13722 41012 13728 41024
rect 13780 41012 13786 41064
rect 13817 41055 13875 41061
rect 13817 41021 13829 41055
rect 13863 41052 13875 41055
rect 14826 41052 14832 41064
rect 13863 41024 14832 41052
rect 13863 41021 13875 41024
rect 13817 41015 13875 41021
rect 14826 41012 14832 41024
rect 14884 41012 14890 41064
rect 14936 41052 14964 41083
rect 15212 41052 15240 41092
rect 17678 41080 17684 41092
rect 17736 41080 17742 41132
rect 18322 41080 18328 41132
rect 18380 41120 18386 41132
rect 22002 41120 22008 41132
rect 18380 41092 22008 41120
rect 18380 41080 18386 41092
rect 22002 41080 22008 41092
rect 22060 41080 22066 41132
rect 19518 41052 19524 41064
rect 14936 41024 15240 41052
rect 19431 41024 19524 41052
rect 19518 41012 19524 41024
rect 19576 41052 19582 41064
rect 19797 41055 19855 41061
rect 19576 41024 19656 41052
rect 19576 41012 19582 41024
rect 12437 40987 12495 40993
rect 12437 40953 12449 40987
rect 12483 40984 12495 40987
rect 13446 40984 13452 40996
rect 12483 40956 13452 40984
rect 12483 40953 12495 40956
rect 12437 40947 12495 40953
rect 12912 40925 12940 40956
rect 13446 40944 13452 40956
rect 13504 40944 13510 40996
rect 16669 40987 16727 40993
rect 16669 40953 16681 40987
rect 16715 40984 16727 40987
rect 17310 40984 17316 40996
rect 16715 40956 17316 40984
rect 16715 40953 16727 40956
rect 16669 40947 16727 40953
rect 17310 40944 17316 40956
rect 17368 40984 17374 40996
rect 17586 40984 17592 40996
rect 17368 40956 17592 40984
rect 17368 40944 17374 40956
rect 17586 40944 17592 40956
rect 17644 40944 17650 40996
rect 19628 40984 19656 41024
rect 19797 41021 19809 41055
rect 19843 41052 19855 41055
rect 20806 41052 20812 41064
rect 19843 41024 20812 41052
rect 19843 41021 19855 41024
rect 19797 41015 19855 41021
rect 20806 41012 20812 41024
rect 20864 41052 20870 41064
rect 21358 41052 21364 41064
rect 20864 41024 21364 41052
rect 20864 41012 20870 41024
rect 21358 41012 21364 41024
rect 21416 41012 21422 41064
rect 21910 41052 21916 41064
rect 21871 41024 21916 41052
rect 21910 41012 21916 41024
rect 21968 41012 21974 41064
rect 20438 40984 20444 40996
rect 19628 40956 20444 40984
rect 20438 40944 20444 40956
rect 20496 40944 20502 40996
rect 23293 40987 23351 40993
rect 23293 40953 23305 40987
rect 23339 40984 23351 40987
rect 23842 40984 23848 40996
rect 23339 40956 23848 40984
rect 23339 40953 23351 40956
rect 23293 40947 23351 40953
rect 12897 40919 12955 40925
rect 12897 40885 12909 40919
rect 12943 40885 12955 40919
rect 13078 40916 13084 40928
rect 13039 40888 13084 40916
rect 12897 40879 12955 40885
rect 13078 40876 13084 40888
rect 13136 40876 13142 40928
rect 13262 40876 13268 40928
rect 13320 40916 13326 40928
rect 15838 40916 15844 40928
rect 13320 40888 15844 40916
rect 13320 40876 13326 40888
rect 15838 40876 15844 40888
rect 15896 40876 15902 40928
rect 15930 40876 15936 40928
rect 15988 40916 15994 40928
rect 16117 40919 16175 40925
rect 15988 40888 16033 40916
rect 15988 40876 15994 40888
rect 16117 40885 16129 40919
rect 16163 40916 16175 40919
rect 17037 40919 17095 40925
rect 17037 40916 17049 40919
rect 16163 40888 17049 40916
rect 16163 40885 16175 40888
rect 16117 40879 16175 40885
rect 17037 40885 17049 40888
rect 17083 40885 17095 40919
rect 17037 40879 17095 40885
rect 18322 40876 18328 40928
rect 18380 40916 18386 40928
rect 19061 40919 19119 40925
rect 19061 40916 19073 40919
rect 18380 40888 19073 40916
rect 18380 40876 18386 40888
rect 19061 40885 19073 40888
rect 19107 40885 19119 40919
rect 19061 40879 19119 40885
rect 21542 40876 21548 40928
rect 21600 40916 21606 40928
rect 23308 40916 23336 40947
rect 23842 40944 23848 40956
rect 23900 40944 23906 40996
rect 21600 40888 23336 40916
rect 21600 40876 21606 40888
rect 1104 40826 38824 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 38824 40826
rect 1104 40752 38824 40774
rect 12250 40712 12256 40724
rect 12211 40684 12256 40712
rect 12250 40672 12256 40684
rect 12308 40672 12314 40724
rect 13078 40712 13084 40724
rect 13039 40684 13084 40712
rect 13078 40672 13084 40684
rect 13136 40672 13142 40724
rect 16298 40672 16304 40724
rect 16356 40712 16362 40724
rect 16853 40715 16911 40721
rect 16853 40712 16865 40715
rect 16356 40684 16865 40712
rect 16356 40672 16362 40684
rect 16853 40681 16865 40684
rect 16899 40681 16911 40715
rect 16853 40675 16911 40681
rect 17034 40672 17040 40724
rect 17092 40712 17098 40724
rect 18049 40715 18107 40721
rect 18049 40712 18061 40715
rect 17092 40684 18061 40712
rect 17092 40672 17098 40684
rect 18049 40681 18061 40684
rect 18095 40681 18107 40715
rect 18049 40675 18107 40681
rect 20625 40715 20683 40721
rect 20625 40681 20637 40715
rect 20671 40712 20683 40715
rect 21450 40712 21456 40724
rect 20671 40684 21456 40712
rect 20671 40681 20683 40684
rect 20625 40675 20683 40681
rect 21450 40672 21456 40684
rect 21508 40672 21514 40724
rect 21634 40672 21640 40724
rect 21692 40712 21698 40724
rect 25406 40712 25412 40724
rect 21692 40684 25412 40712
rect 21692 40672 21698 40684
rect 25406 40672 25412 40684
rect 25464 40672 25470 40724
rect 12161 40647 12219 40653
rect 12161 40613 12173 40647
rect 12207 40644 12219 40647
rect 12207 40616 12434 40644
rect 12207 40613 12219 40616
rect 12161 40607 12219 40613
rect 12406 40508 12434 40616
rect 16390 40604 16396 40656
rect 16448 40644 16454 40656
rect 19518 40644 19524 40656
rect 16448 40616 19524 40644
rect 16448 40604 16454 40616
rect 19518 40604 19524 40616
rect 19576 40604 19582 40656
rect 14642 40576 14648 40588
rect 14603 40548 14648 40576
rect 14642 40536 14648 40548
rect 14700 40536 14706 40588
rect 16942 40576 16948 40588
rect 16040 40548 16948 40576
rect 12526 40508 12532 40520
rect 12406 40480 12532 40508
rect 12526 40468 12532 40480
rect 12584 40508 12590 40520
rect 12713 40511 12771 40517
rect 12713 40508 12725 40511
rect 12584 40480 12725 40508
rect 12584 40468 12590 40480
rect 12713 40477 12725 40480
rect 12759 40477 12771 40511
rect 14660 40508 14688 40536
rect 15930 40508 15936 40520
rect 14660 40480 15936 40508
rect 12713 40471 12771 40477
rect 15930 40468 15936 40480
rect 15988 40468 15994 40520
rect 11793 40443 11851 40449
rect 11793 40409 11805 40443
rect 11839 40440 11851 40443
rect 13170 40440 13176 40452
rect 11839 40412 13176 40440
rect 11839 40409 11851 40412
rect 11793 40403 11851 40409
rect 13170 40400 13176 40412
rect 13228 40400 13234 40452
rect 14918 40449 14924 40452
rect 14912 40403 14924 40449
rect 14976 40440 14982 40452
rect 14976 40412 15012 40440
rect 14918 40400 14924 40403
rect 14976 40400 14982 40412
rect 13078 40372 13084 40384
rect 13039 40344 13084 40372
rect 13078 40332 13084 40344
rect 13136 40332 13142 40384
rect 13262 40372 13268 40384
rect 13223 40344 13268 40372
rect 13262 40332 13268 40344
rect 13320 40332 13326 40384
rect 16040 40381 16068 40548
rect 16942 40536 16948 40548
rect 17000 40576 17006 40588
rect 21174 40576 21180 40588
rect 17000 40548 18184 40576
rect 17000 40536 17006 40548
rect 16482 40508 16488 40520
rect 16443 40480 16488 40508
rect 16482 40468 16488 40480
rect 16540 40468 16546 40520
rect 16669 40511 16727 40517
rect 16669 40508 16681 40511
rect 16592 40480 16681 40508
rect 16592 40384 16620 40480
rect 16669 40477 16681 40480
rect 16715 40508 16727 40511
rect 16758 40508 16764 40520
rect 16715 40480 16764 40508
rect 16715 40477 16727 40480
rect 16669 40471 16727 40477
rect 16758 40468 16764 40480
rect 16816 40468 16822 40520
rect 17310 40508 17316 40520
rect 17271 40480 17316 40508
rect 17310 40468 17316 40480
rect 17368 40468 17374 40520
rect 17506 40517 17534 40548
rect 17497 40511 17555 40517
rect 17497 40477 17509 40511
rect 17543 40477 17555 40511
rect 17954 40508 17960 40520
rect 17915 40480 17960 40508
rect 17497 40471 17555 40477
rect 17954 40468 17960 40480
rect 18012 40468 18018 40520
rect 18156 40517 18184 40548
rect 21008 40548 21180 40576
rect 18141 40511 18199 40517
rect 18141 40477 18153 40511
rect 18187 40477 18199 40511
rect 18141 40471 18199 40477
rect 19334 40468 19340 40520
rect 19392 40508 19398 40520
rect 19613 40511 19671 40517
rect 19613 40508 19625 40511
rect 19392 40480 19625 40508
rect 19392 40468 19398 40480
rect 19613 40477 19625 40480
rect 19659 40477 19671 40511
rect 19613 40471 19671 40477
rect 20806 40468 20812 40520
rect 20864 40517 20870 40520
rect 21008 40517 21036 40548
rect 21174 40536 21180 40548
rect 21232 40576 21238 40588
rect 21232 40548 22232 40576
rect 21232 40536 21238 40548
rect 20864 40511 20913 40517
rect 20864 40477 20867 40511
rect 20901 40477 20913 40511
rect 20864 40471 20913 40477
rect 20990 40511 21048 40517
rect 20990 40477 21002 40511
rect 21036 40477 21048 40511
rect 20990 40471 21048 40477
rect 21085 40511 21143 40517
rect 21085 40477 21097 40511
rect 21131 40477 21143 40511
rect 21085 40471 21143 40477
rect 21269 40511 21327 40517
rect 21269 40477 21281 40511
rect 21315 40508 21327 40511
rect 21358 40508 21364 40520
rect 21315 40480 21364 40508
rect 21315 40477 21327 40480
rect 21269 40471 21327 40477
rect 20864 40468 20870 40471
rect 21100 40456 21133 40471
rect 21358 40468 21364 40480
rect 21416 40508 21422 40520
rect 21416 40480 21956 40508
rect 21416 40468 21422 40480
rect 17405 40443 17463 40449
rect 17405 40409 17417 40443
rect 17451 40440 17463 40443
rect 17586 40440 17592 40452
rect 17451 40412 17592 40440
rect 17451 40409 17463 40412
rect 17405 40403 17463 40409
rect 17586 40400 17592 40412
rect 17644 40400 17650 40452
rect 21105 40440 21133 40456
rect 21818 40440 21824 40452
rect 21105 40412 21189 40440
rect 21779 40412 21824 40440
rect 16025 40375 16083 40381
rect 16025 40341 16037 40375
rect 16071 40341 16083 40375
rect 16025 40335 16083 40341
rect 16574 40332 16580 40384
rect 16632 40332 16638 40384
rect 16850 40332 16856 40384
rect 16908 40372 16914 40384
rect 17218 40372 17224 40384
rect 16908 40344 17224 40372
rect 16908 40332 16914 40344
rect 17218 40332 17224 40344
rect 17276 40372 17282 40384
rect 18782 40372 18788 40384
rect 17276 40344 18788 40372
rect 17276 40332 17282 40344
rect 18782 40332 18788 40344
rect 18840 40332 18846 40384
rect 19429 40375 19487 40381
rect 19429 40341 19441 40375
rect 19475 40372 19487 40375
rect 20254 40372 20260 40384
rect 19475 40344 20260 40372
rect 19475 40341 19487 40344
rect 19429 40335 19487 40341
rect 20254 40332 20260 40344
rect 20312 40332 20318 40384
rect 21161 40372 21189 40412
rect 21818 40400 21824 40412
rect 21876 40400 21882 40452
rect 21928 40440 21956 40480
rect 22002 40468 22008 40520
rect 22060 40508 22066 40520
rect 22204 40517 22232 40548
rect 22097 40511 22155 40517
rect 22097 40508 22109 40511
rect 22060 40480 22109 40508
rect 22060 40468 22066 40480
rect 22097 40477 22109 40480
rect 22143 40477 22155 40511
rect 22097 40471 22155 40477
rect 22189 40511 22247 40517
rect 22189 40477 22201 40511
rect 22235 40477 22247 40511
rect 22189 40471 22247 40477
rect 22278 40468 22284 40520
rect 22336 40517 22342 40520
rect 22336 40508 22344 40517
rect 22465 40511 22523 40517
rect 22336 40480 22381 40508
rect 22336 40471 22344 40480
rect 22465 40477 22477 40511
rect 22511 40477 22523 40511
rect 22465 40471 22523 40477
rect 22336 40468 22342 40471
rect 22480 40440 22508 40471
rect 21928 40412 22508 40440
rect 22830 40372 22836 40384
rect 21161 40344 22836 40372
rect 22830 40332 22836 40344
rect 22888 40332 22894 40384
rect 1104 40282 38824 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 38824 40282
rect 1104 40208 38824 40230
rect 17862 40168 17868 40180
rect 15488 40140 17868 40168
rect 13262 40060 13268 40112
rect 13320 40100 13326 40112
rect 15488 40109 15516 40140
rect 17862 40128 17868 40140
rect 17920 40128 17926 40180
rect 19242 40168 19248 40180
rect 19203 40140 19248 40168
rect 19242 40128 19248 40140
rect 19300 40128 19306 40180
rect 19904 40140 22600 40168
rect 15473 40103 15531 40109
rect 13320 40072 14872 40100
rect 13320 40060 13326 40072
rect 11793 40035 11851 40041
rect 11793 40001 11805 40035
rect 11839 40032 11851 40035
rect 12066 40032 12072 40044
rect 11839 40004 12072 40032
rect 11839 40001 11851 40004
rect 11793 39995 11851 40001
rect 12066 39992 12072 40004
rect 12124 39992 12130 40044
rect 12805 40035 12863 40041
rect 12805 40001 12817 40035
rect 12851 40032 12863 40035
rect 12894 40032 12900 40044
rect 12851 40004 12900 40032
rect 12851 40001 12863 40004
rect 12805 39995 12863 40001
rect 12894 39992 12900 40004
rect 12952 39992 12958 40044
rect 14844 40041 14872 40072
rect 15473 40069 15485 40103
rect 15519 40069 15531 40103
rect 15473 40063 15531 40069
rect 15657 40103 15715 40109
rect 15657 40069 15669 40103
rect 15703 40100 15715 40103
rect 16942 40100 16948 40112
rect 15703 40072 16948 40100
rect 15703 40069 15715 40072
rect 15657 40063 15715 40069
rect 16942 40060 16948 40072
rect 17000 40060 17006 40112
rect 19904 40109 19932 40140
rect 19889 40103 19947 40109
rect 19889 40069 19901 40103
rect 19935 40069 19947 40103
rect 20089 40103 20147 40109
rect 20089 40100 20101 40103
rect 19889 40063 19947 40069
rect 19996 40072 20101 40100
rect 13072 40035 13130 40041
rect 13072 40001 13084 40035
rect 13118 40032 13130 40035
rect 14829 40035 14887 40041
rect 13118 40004 14688 40032
rect 13118 40001 13130 40004
rect 13072 39995 13130 40001
rect 11514 39964 11520 39976
rect 11475 39936 11520 39964
rect 11514 39924 11520 39936
rect 11572 39924 11578 39976
rect 14660 39905 14688 40004
rect 14829 40001 14841 40035
rect 14875 40001 14887 40035
rect 14829 39995 14887 40001
rect 17218 39992 17224 40044
rect 17276 40032 17282 40044
rect 18325 40035 18383 40041
rect 18325 40032 18337 40035
rect 17276 40004 18337 40032
rect 17276 39992 17282 40004
rect 18325 40001 18337 40004
rect 18371 40001 18383 40035
rect 18506 40032 18512 40044
rect 18467 40004 18512 40032
rect 18325 39995 18383 40001
rect 18506 39992 18512 40004
rect 18564 39992 18570 40044
rect 18785 40035 18843 40041
rect 18785 40001 18797 40035
rect 18831 40032 18843 40035
rect 19996 40032 20024 40072
rect 20089 40069 20101 40072
rect 20135 40069 20147 40103
rect 20089 40063 20147 40069
rect 20254 40060 20260 40112
rect 20312 40100 20318 40112
rect 20901 40103 20959 40109
rect 20901 40100 20913 40103
rect 20312 40072 20913 40100
rect 20312 40060 20318 40072
rect 20901 40069 20913 40072
rect 20947 40069 20959 40103
rect 20901 40063 20959 40069
rect 21085 40103 21143 40109
rect 21085 40069 21097 40103
rect 21131 40100 21143 40103
rect 21542 40100 21548 40112
rect 21131 40072 21548 40100
rect 21131 40069 21143 40072
rect 21085 40063 21143 40069
rect 21542 40060 21548 40072
rect 21600 40060 21606 40112
rect 22572 40100 22600 40140
rect 23198 40128 23204 40180
rect 23256 40168 23262 40180
rect 24137 40171 24195 40177
rect 24137 40168 24149 40171
rect 23256 40140 24149 40168
rect 23256 40128 23262 40140
rect 24137 40137 24149 40140
rect 24183 40137 24195 40171
rect 24137 40131 24195 40137
rect 23937 40103 23995 40109
rect 23937 40100 23949 40103
rect 22572 40072 23949 40100
rect 23937 40069 23949 40072
rect 23983 40100 23995 40103
rect 25498 40100 25504 40112
rect 23983 40072 25504 40100
rect 23983 40069 23995 40072
rect 23937 40063 23995 40069
rect 25498 40060 25504 40072
rect 25556 40060 25562 40112
rect 18831 40004 20024 40032
rect 21269 40035 21327 40041
rect 18831 40001 18843 40004
rect 18785 39995 18843 40001
rect 21269 40001 21281 40035
rect 21315 40032 21327 40035
rect 22278 40032 22284 40044
rect 21315 40004 22284 40032
rect 21315 40001 21327 40004
rect 21269 39995 21327 40001
rect 15102 39924 15108 39976
rect 15160 39964 15166 39976
rect 17310 39964 17316 39976
rect 15160 39936 17316 39964
rect 15160 39924 15166 39936
rect 17310 39924 17316 39936
rect 17368 39964 17374 39976
rect 17954 39964 17960 39976
rect 17368 39936 17960 39964
rect 17368 39924 17374 39936
rect 17954 39924 17960 39936
rect 18012 39924 18018 39976
rect 18417 39967 18475 39973
rect 18417 39933 18429 39967
rect 18463 39964 18475 39967
rect 18800 39964 18828 39995
rect 22278 39992 22284 40004
rect 22336 39992 22342 40044
rect 24854 40032 24860 40044
rect 24815 40004 24860 40032
rect 24854 39992 24860 40004
rect 24912 39992 24918 40044
rect 25038 40032 25044 40044
rect 24999 40004 25044 40032
rect 25038 39992 25044 40004
rect 25096 39992 25102 40044
rect 18463 39936 18828 39964
rect 23017 39967 23075 39973
rect 18463 39933 18475 39936
rect 18417 39927 18475 39933
rect 23017 39933 23029 39967
rect 23063 39964 23075 39967
rect 23198 39964 23204 39976
rect 23063 39936 23204 39964
rect 23063 39933 23075 39936
rect 23017 39927 23075 39933
rect 23198 39924 23204 39936
rect 23256 39924 23262 39976
rect 14645 39899 14703 39905
rect 14645 39865 14657 39899
rect 14691 39865 14703 39899
rect 14645 39859 14703 39865
rect 15654 39856 15660 39908
rect 15712 39896 15718 39908
rect 16298 39896 16304 39908
rect 15712 39868 16304 39896
rect 15712 39856 15718 39868
rect 16298 39856 16304 39868
rect 16356 39856 16362 39908
rect 19153 39899 19211 39905
rect 19153 39865 19165 39899
rect 19199 39896 19211 39899
rect 19334 39896 19340 39908
rect 19199 39868 19340 39896
rect 19199 39865 19211 39868
rect 19153 39859 19211 39865
rect 19334 39856 19340 39868
rect 19392 39856 19398 39908
rect 19613 39899 19671 39905
rect 19613 39865 19625 39899
rect 19659 39896 19671 39899
rect 20530 39896 20536 39908
rect 19659 39868 20536 39896
rect 19659 39865 19671 39868
rect 19613 39859 19671 39865
rect 14182 39828 14188 39840
rect 14143 39800 14188 39828
rect 14182 39788 14188 39800
rect 14240 39788 14246 39840
rect 15378 39788 15384 39840
rect 15436 39828 15442 39840
rect 20088 39837 20116 39868
rect 20530 39856 20536 39868
rect 20588 39856 20594 39908
rect 23290 39896 23296 39908
rect 23251 39868 23296 39896
rect 23290 39856 23296 39868
rect 23348 39856 23354 39908
rect 23474 39896 23480 39908
rect 23435 39868 23480 39896
rect 23474 39856 23480 39868
rect 23532 39856 23538 39908
rect 24136 39868 31754 39896
rect 15841 39831 15899 39837
rect 15841 39828 15853 39831
rect 15436 39800 15853 39828
rect 15436 39788 15442 39800
rect 15841 39797 15853 39800
rect 15887 39797 15899 39831
rect 15841 39791 15899 39797
rect 20073 39831 20131 39837
rect 20073 39797 20085 39831
rect 20119 39797 20131 39831
rect 20254 39828 20260 39840
rect 20215 39800 20260 39828
rect 20073 39791 20131 39797
rect 20254 39788 20260 39800
rect 20312 39788 20318 39840
rect 24136 39837 24164 39868
rect 24121 39831 24179 39837
rect 24121 39797 24133 39831
rect 24167 39797 24179 39831
rect 24302 39828 24308 39840
rect 24263 39800 24308 39828
rect 24121 39791 24179 39797
rect 24302 39788 24308 39800
rect 24360 39788 24366 39840
rect 31726 39828 31754 39868
rect 36170 39828 36176 39840
rect 31726 39800 36176 39828
rect 36170 39788 36176 39800
rect 36228 39788 36234 39840
rect 1104 39738 38824 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 38824 39738
rect 1104 39664 38824 39686
rect 12526 39624 12532 39636
rect 12487 39596 12532 39624
rect 12526 39584 12532 39596
rect 12584 39584 12590 39636
rect 13078 39584 13084 39636
rect 13136 39624 13142 39636
rect 13265 39627 13323 39633
rect 13265 39624 13277 39627
rect 13136 39596 13277 39624
rect 13136 39584 13142 39596
rect 13265 39593 13277 39596
rect 13311 39593 13323 39627
rect 14918 39624 14924 39636
rect 14879 39596 14924 39624
rect 13265 39587 13323 39593
rect 14918 39584 14924 39596
rect 14976 39584 14982 39636
rect 16758 39624 16764 39636
rect 15028 39596 16764 39624
rect 12636 39460 13216 39488
rect 12636 39432 12664 39460
rect 11609 39423 11667 39429
rect 11609 39389 11621 39423
rect 11655 39420 11667 39423
rect 12250 39420 12256 39432
rect 11655 39392 12256 39420
rect 11655 39389 11667 39392
rect 11609 39383 11667 39389
rect 12250 39380 12256 39392
rect 12308 39380 12314 39432
rect 12529 39423 12587 39429
rect 12529 39389 12541 39423
rect 12575 39420 12587 39423
rect 12618 39420 12624 39432
rect 12575 39392 12624 39420
rect 12575 39389 12587 39392
rect 12529 39383 12587 39389
rect 12618 39380 12624 39392
rect 12676 39380 12682 39432
rect 13188 39429 13216 39460
rect 12713 39423 12771 39429
rect 12713 39389 12725 39423
rect 12759 39389 12771 39423
rect 12713 39383 12771 39389
rect 13173 39423 13231 39429
rect 13173 39389 13185 39423
rect 13219 39389 13231 39423
rect 13173 39383 13231 39389
rect 13357 39423 13415 39429
rect 13357 39389 13369 39423
rect 13403 39420 13415 39423
rect 15028 39420 15056 39596
rect 16758 39584 16764 39596
rect 16816 39584 16822 39636
rect 24854 39584 24860 39636
rect 24912 39624 24918 39636
rect 25225 39627 25283 39633
rect 25225 39624 25237 39627
rect 24912 39596 25237 39624
rect 24912 39584 24918 39596
rect 25225 39593 25237 39596
rect 25271 39593 25283 39627
rect 25225 39587 25283 39593
rect 25406 39584 25412 39636
rect 25464 39624 25470 39636
rect 25501 39627 25559 39633
rect 25501 39624 25513 39627
rect 25464 39596 25513 39624
rect 25464 39584 25470 39596
rect 25501 39593 25513 39596
rect 25547 39593 25559 39627
rect 25501 39587 25559 39593
rect 26053 39627 26111 39633
rect 26053 39593 26065 39627
rect 26099 39624 26111 39627
rect 32950 39624 32956 39636
rect 26099 39596 32956 39624
rect 26099 39593 26111 39596
rect 26053 39587 26111 39593
rect 25130 39556 25136 39568
rect 25091 39528 25136 39556
rect 25130 39516 25136 39528
rect 25188 39516 25194 39568
rect 15654 39488 15660 39500
rect 15304 39460 15660 39488
rect 15304 39429 15332 39460
rect 15654 39448 15660 39460
rect 15712 39448 15718 39500
rect 15930 39448 15936 39500
rect 15988 39488 15994 39500
rect 16025 39491 16083 39497
rect 16025 39488 16037 39491
rect 15988 39460 16037 39488
rect 15988 39448 15994 39460
rect 16025 39457 16037 39460
rect 16071 39457 16083 39491
rect 16025 39451 16083 39457
rect 13403 39392 15056 39420
rect 15197 39423 15255 39429
rect 13403 39389 13415 39392
rect 13357 39383 13415 39389
rect 15197 39389 15209 39423
rect 15243 39389 15255 39423
rect 15197 39383 15255 39389
rect 15289 39423 15347 39429
rect 15289 39389 15301 39423
rect 15335 39389 15347 39423
rect 15289 39383 15347 39389
rect 12728 39352 12756 39383
rect 13372 39352 13400 39383
rect 12728 39324 13400 39352
rect 14274 39312 14280 39364
rect 14332 39352 14338 39364
rect 15212 39352 15240 39383
rect 15378 39380 15384 39432
rect 15436 39420 15442 39432
rect 15565 39423 15623 39429
rect 15436 39392 15481 39420
rect 15436 39380 15442 39392
rect 15565 39389 15577 39423
rect 15611 39420 15623 39423
rect 15838 39420 15844 39432
rect 15611 39392 15844 39420
rect 15611 39389 15623 39392
rect 15565 39383 15623 39389
rect 15838 39380 15844 39392
rect 15896 39380 15902 39432
rect 19426 39420 19432 39432
rect 19387 39392 19432 39420
rect 19426 39380 19432 39392
rect 19484 39380 19490 39432
rect 19889 39423 19947 39429
rect 19889 39389 19901 39423
rect 19935 39420 19947 39423
rect 21082 39420 21088 39432
rect 19935 39392 21088 39420
rect 19935 39389 19947 39392
rect 19889 39383 19947 39389
rect 21082 39380 21088 39392
rect 21140 39380 21146 39432
rect 21910 39420 21916 39432
rect 21871 39392 21916 39420
rect 21910 39380 21916 39392
rect 21968 39380 21974 39432
rect 25516 39420 25544 39587
rect 32950 39584 32956 39596
rect 33008 39584 33014 39636
rect 25516 39392 25912 39420
rect 14332 39324 15332 39352
rect 14332 39312 14338 39324
rect 15304 39296 15332 39324
rect 15470 39312 15476 39364
rect 15528 39352 15534 39364
rect 16270 39355 16328 39361
rect 16270 39352 16282 39355
rect 15528 39324 16282 39352
rect 15528 39312 15534 39324
rect 16270 39321 16282 39324
rect 16316 39321 16328 39355
rect 17862 39352 17868 39364
rect 17823 39324 17868 39352
rect 16270 39315 16328 39321
rect 17862 39312 17868 39324
rect 17920 39312 17926 39364
rect 18049 39355 18107 39361
rect 18049 39321 18061 39355
rect 18095 39352 18107 39355
rect 18506 39352 18512 39364
rect 18095 39324 18512 39352
rect 18095 39321 18107 39324
rect 18049 39315 18107 39321
rect 18506 39312 18512 39324
rect 18564 39312 18570 39364
rect 20990 39352 20996 39364
rect 20951 39324 20996 39352
rect 20990 39312 20996 39324
rect 21048 39312 21054 39364
rect 22186 39361 22192 39364
rect 21177 39355 21235 39361
rect 21177 39321 21189 39355
rect 21223 39352 21235 39355
rect 21223 39324 22094 39352
rect 21223 39321 21235 39324
rect 21177 39315 21235 39321
rect 22066 39296 22094 39324
rect 22180 39315 22192 39361
rect 22244 39352 22250 39364
rect 24765 39355 24823 39361
rect 22244 39324 22280 39352
rect 22186 39312 22192 39315
rect 22244 39312 22250 39324
rect 24765 39321 24777 39355
rect 24811 39352 24823 39355
rect 24854 39352 24860 39364
rect 24811 39324 24860 39352
rect 24811 39321 24823 39324
rect 24765 39315 24823 39321
rect 24854 39312 24860 39324
rect 24912 39352 24918 39364
rect 25884 39361 25912 39392
rect 25869 39355 25927 39361
rect 24912 39324 25636 39352
rect 24912 39312 24918 39324
rect 11425 39287 11483 39293
rect 11425 39253 11437 39287
rect 11471 39284 11483 39287
rect 11606 39284 11612 39296
rect 11471 39256 11612 39284
rect 11471 39253 11483 39256
rect 11425 39247 11483 39253
rect 11606 39244 11612 39256
rect 11664 39244 11670 39296
rect 15286 39244 15292 39296
rect 15344 39244 15350 39296
rect 17218 39244 17224 39296
rect 17276 39284 17282 39296
rect 17405 39287 17463 39293
rect 17405 39284 17417 39287
rect 17276 39256 17417 39284
rect 17276 39244 17282 39256
rect 17405 39253 17417 39256
rect 17451 39253 17463 39287
rect 18230 39284 18236 39296
rect 18191 39256 18236 39284
rect 17405 39247 17463 39253
rect 18230 39244 18236 39256
rect 18288 39244 18294 39296
rect 19245 39287 19303 39293
rect 19245 39253 19257 39287
rect 19291 39284 19303 39287
rect 20070 39284 20076 39296
rect 19291 39256 20076 39284
rect 19291 39253 19303 39256
rect 19245 39247 19303 39253
rect 20070 39244 20076 39256
rect 20128 39244 20134 39296
rect 20530 39284 20536 39296
rect 20491 39256 20536 39284
rect 20530 39244 20536 39256
rect 20588 39244 20594 39296
rect 21361 39287 21419 39293
rect 21361 39253 21373 39287
rect 21407 39284 21419 39287
rect 21450 39284 21456 39296
rect 21407 39256 21456 39284
rect 21407 39253 21419 39256
rect 21361 39247 21419 39253
rect 21450 39244 21456 39256
rect 21508 39244 21514 39296
rect 22066 39256 22100 39296
rect 22094 39244 22100 39256
rect 22152 39284 22158 39296
rect 23293 39287 23351 39293
rect 23293 39284 23305 39287
rect 22152 39256 23305 39284
rect 22152 39244 22158 39256
rect 23293 39253 23305 39256
rect 23339 39253 23351 39287
rect 25608 39284 25636 39324
rect 25869 39321 25881 39355
rect 25915 39352 25927 39355
rect 25958 39352 25964 39364
rect 25915 39324 25964 39352
rect 25915 39321 25927 39324
rect 25869 39315 25927 39321
rect 25958 39312 25964 39324
rect 26016 39312 26022 39364
rect 26069 39287 26127 39293
rect 26069 39284 26081 39287
rect 25608 39256 26081 39284
rect 23293 39247 23351 39253
rect 26069 39253 26081 39256
rect 26115 39253 26127 39287
rect 26234 39284 26240 39296
rect 26195 39256 26240 39284
rect 26069 39247 26127 39253
rect 26234 39244 26240 39256
rect 26292 39244 26298 39296
rect 1104 39194 38824 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 38824 39194
rect 1104 39120 38824 39142
rect 11514 39040 11520 39092
rect 11572 39080 11578 39092
rect 12069 39083 12127 39089
rect 12069 39080 12081 39083
rect 11572 39052 12081 39080
rect 11572 39040 11578 39052
rect 12069 39049 12081 39052
rect 12115 39049 12127 39083
rect 15470 39080 15476 39092
rect 15431 39052 15476 39080
rect 12069 39043 12127 39049
rect 15470 39040 15476 39052
rect 15528 39040 15534 39092
rect 15930 39040 15936 39092
rect 15988 39080 15994 39092
rect 15988 39052 17540 39080
rect 15988 39040 15994 39052
rect 15654 38972 15660 39024
rect 15712 39012 15718 39024
rect 17310 39012 17316 39024
rect 15712 38984 17316 39012
rect 15712 38972 15718 38984
rect 15856 38953 15884 38984
rect 17310 38972 17316 38984
rect 17368 38972 17374 39024
rect 15749 38947 15807 38953
rect 15749 38913 15761 38947
rect 15795 38913 15807 38947
rect 15749 38907 15807 38913
rect 15841 38947 15899 38953
rect 15841 38913 15853 38947
rect 15887 38913 15899 38947
rect 15841 38907 15899 38913
rect 11609 38879 11667 38885
rect 11609 38845 11621 38879
rect 11655 38876 11667 38879
rect 12526 38876 12532 38888
rect 11655 38848 12532 38876
rect 11655 38845 11667 38848
rect 11609 38839 11667 38845
rect 12526 38836 12532 38848
rect 12584 38836 12590 38888
rect 15764 38876 15792 38907
rect 15930 38904 15936 38956
rect 15988 38944 15994 38956
rect 17512 38953 17540 39052
rect 21082 39040 21088 39092
rect 21140 39080 21146 39092
rect 21177 39083 21235 39089
rect 21177 39080 21189 39083
rect 21140 39052 21189 39080
rect 21140 39040 21146 39052
rect 21177 39049 21189 39052
rect 21223 39049 21235 39083
rect 21177 39043 21235 39049
rect 26237 39083 26295 39089
rect 26237 39049 26249 39083
rect 26283 39049 26295 39083
rect 26237 39043 26295 39049
rect 21910 39012 21916 39024
rect 19812 38984 21916 39012
rect 16117 38947 16175 38953
rect 15988 38916 16033 38944
rect 15988 38904 15994 38916
rect 16117 38913 16129 38947
rect 16163 38944 16175 38947
rect 17497 38947 17555 38953
rect 16163 38916 17356 38944
rect 16163 38913 16175 38916
rect 16117 38907 16175 38913
rect 16022 38876 16028 38888
rect 15764 38848 16028 38876
rect 16022 38836 16028 38848
rect 16080 38876 16086 38888
rect 16390 38876 16396 38888
rect 16080 38848 16396 38876
rect 16080 38836 16086 38848
rect 16390 38836 16396 38848
rect 16448 38836 16454 38888
rect 11882 38808 11888 38820
rect 11843 38780 11888 38808
rect 11882 38768 11888 38780
rect 11940 38768 11946 38820
rect 17328 38740 17356 38916
rect 17497 38913 17509 38947
rect 17543 38913 17555 38947
rect 17497 38907 17555 38913
rect 17586 38904 17592 38956
rect 17644 38944 17650 38956
rect 19812 38953 19840 38984
rect 21910 38972 21916 38984
rect 21968 39012 21974 39024
rect 21968 38984 22094 39012
rect 21968 38972 21974 38984
rect 20070 38953 20076 38956
rect 17753 38947 17811 38953
rect 17753 38944 17765 38947
rect 17644 38916 17765 38944
rect 17644 38904 17650 38916
rect 17753 38913 17765 38916
rect 17799 38913 17811 38947
rect 17753 38907 17811 38913
rect 19797 38947 19855 38953
rect 19797 38913 19809 38947
rect 19843 38913 19855 38947
rect 20064 38944 20076 38953
rect 20031 38916 20076 38944
rect 19797 38907 19855 38913
rect 20064 38907 20076 38916
rect 20070 38904 20076 38907
rect 20128 38904 20134 38956
rect 22066 38944 22094 38984
rect 22278 38972 22284 39024
rect 22336 39012 22342 39024
rect 22618 39015 22676 39021
rect 22618 39012 22630 39015
rect 22336 38984 22630 39012
rect 22336 38972 22342 38984
rect 22618 38981 22630 38984
rect 22664 38981 22676 39015
rect 22618 38975 22676 38981
rect 24664 39015 24722 39021
rect 24664 38981 24676 39015
rect 24710 39012 24722 39015
rect 26252 39012 26280 39043
rect 24710 38984 26280 39012
rect 24710 38981 24722 38984
rect 24664 38975 24722 38981
rect 22373 38947 22431 38953
rect 22373 38944 22385 38947
rect 22066 38916 22385 38944
rect 22373 38913 22385 38916
rect 22419 38913 22431 38947
rect 26418 38944 26424 38956
rect 26379 38916 26424 38944
rect 22373 38907 22431 38913
rect 26418 38904 26424 38916
rect 26476 38904 26482 38956
rect 24397 38879 24455 38885
rect 24397 38845 24409 38879
rect 24443 38845 24455 38879
rect 24397 38839 24455 38845
rect 17678 38740 17684 38752
rect 17328 38712 17684 38740
rect 17678 38700 17684 38712
rect 17736 38700 17742 38752
rect 18506 38700 18512 38752
rect 18564 38740 18570 38752
rect 18877 38743 18935 38749
rect 18877 38740 18889 38743
rect 18564 38712 18889 38740
rect 18564 38700 18570 38712
rect 18877 38709 18889 38712
rect 18923 38709 18935 38743
rect 23750 38740 23756 38752
rect 23711 38712 23756 38740
rect 18877 38703 18935 38709
rect 23750 38700 23756 38712
rect 23808 38700 23814 38752
rect 24412 38740 24440 38839
rect 25038 38740 25044 38752
rect 24412 38712 25044 38740
rect 25038 38700 25044 38712
rect 25096 38700 25102 38752
rect 25314 38700 25320 38752
rect 25372 38740 25378 38752
rect 25777 38743 25835 38749
rect 25777 38740 25789 38743
rect 25372 38712 25789 38740
rect 25372 38700 25378 38712
rect 25777 38709 25789 38712
rect 25823 38709 25835 38743
rect 25777 38703 25835 38709
rect 1104 38650 38824 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 38824 38650
rect 1104 38576 38824 38598
rect 12710 38536 12716 38548
rect 12671 38508 12716 38536
rect 12710 38496 12716 38508
rect 12768 38536 12774 38548
rect 13265 38539 13323 38545
rect 13265 38536 13277 38539
rect 12768 38508 13277 38536
rect 12768 38496 12774 38508
rect 13265 38505 13277 38508
rect 13311 38505 13323 38539
rect 13265 38499 13323 38505
rect 15841 38539 15899 38545
rect 15841 38505 15853 38539
rect 15887 38536 15899 38539
rect 15930 38536 15936 38548
rect 15887 38508 15936 38536
rect 15887 38505 15899 38508
rect 15841 38499 15899 38505
rect 15930 38496 15936 38508
rect 15988 38496 15994 38548
rect 17218 38536 17224 38548
rect 16224 38508 17224 38536
rect 16224 38468 16252 38508
rect 17218 38496 17224 38508
rect 17276 38496 17282 38548
rect 17313 38539 17371 38545
rect 17313 38505 17325 38539
rect 17359 38536 17371 38539
rect 17586 38536 17592 38548
rect 17359 38508 17592 38536
rect 17359 38505 17371 38508
rect 17313 38499 17371 38505
rect 17586 38496 17592 38508
rect 17644 38496 17650 38548
rect 17678 38496 17684 38548
rect 17736 38536 17742 38548
rect 18046 38536 18052 38548
rect 17736 38508 18052 38536
rect 17736 38496 17742 38508
rect 18046 38496 18052 38508
rect 18104 38496 18110 38548
rect 19797 38539 19855 38545
rect 19797 38505 19809 38539
rect 19843 38536 19855 38539
rect 20254 38536 20260 38548
rect 19843 38508 20260 38536
rect 19843 38505 19855 38508
rect 19797 38499 19855 38505
rect 20254 38496 20260 38508
rect 20312 38496 20318 38548
rect 20806 38496 20812 38548
rect 20864 38536 20870 38548
rect 21174 38536 21180 38548
rect 20864 38508 21180 38536
rect 20864 38496 20870 38508
rect 21174 38496 21180 38508
rect 21232 38496 21238 38548
rect 22097 38539 22155 38545
rect 22097 38505 22109 38539
rect 22143 38536 22155 38539
rect 22278 38536 22284 38548
rect 22143 38508 22284 38536
rect 22143 38505 22155 38508
rect 22097 38499 22155 38505
rect 22278 38496 22284 38508
rect 22336 38496 22342 38548
rect 23198 38536 23204 38548
rect 23159 38508 23204 38536
rect 23198 38496 23204 38508
rect 23256 38496 23262 38548
rect 25501 38539 25559 38545
rect 25501 38505 25513 38539
rect 25547 38536 25559 38539
rect 26234 38536 26240 38548
rect 25547 38508 26240 38536
rect 25547 38505 25559 38508
rect 25501 38499 25559 38505
rect 26234 38496 26240 38508
rect 26292 38496 26298 38548
rect 15672 38440 16252 38468
rect 16316 38440 18368 38468
rect 12345 38403 12403 38409
rect 12345 38369 12357 38403
rect 12391 38400 12403 38403
rect 12434 38400 12440 38412
rect 12391 38372 12440 38400
rect 12391 38369 12403 38372
rect 12345 38363 12403 38369
rect 12434 38360 12440 38372
rect 12492 38400 12498 38412
rect 12894 38400 12900 38412
rect 12492 38372 12900 38400
rect 12492 38360 12498 38372
rect 12894 38360 12900 38372
rect 12952 38360 12958 38412
rect 15194 38400 15200 38412
rect 14200 38372 15200 38400
rect 10689 38335 10747 38341
rect 10689 38301 10701 38335
rect 10735 38332 10747 38335
rect 14200 38332 14228 38372
rect 15194 38360 15200 38372
rect 15252 38360 15258 38412
rect 10735 38304 14228 38332
rect 10735 38301 10747 38304
rect 10689 38295 10747 38301
rect 14274 38292 14280 38344
rect 14332 38332 14338 38344
rect 14332 38304 14377 38332
rect 14332 38292 14338 38304
rect 14918 38292 14924 38344
rect 14976 38332 14982 38344
rect 15672 38341 15700 38440
rect 16316 38341 16344 38440
rect 16850 38400 16856 38412
rect 16592 38372 16856 38400
rect 16592 38341 16620 38372
rect 16850 38360 16856 38372
rect 16908 38360 16914 38412
rect 17310 38360 17316 38412
rect 17368 38400 17374 38412
rect 18230 38400 18236 38412
rect 17368 38372 17724 38400
rect 17368 38360 17374 38372
rect 15657 38335 15715 38341
rect 15657 38332 15669 38335
rect 14976 38304 15669 38332
rect 14976 38292 14982 38304
rect 15657 38301 15669 38304
rect 15703 38301 15715 38335
rect 15657 38295 15715 38301
rect 16301 38335 16359 38341
rect 16301 38301 16313 38335
rect 16347 38301 16359 38335
rect 16301 38295 16359 38301
rect 16577 38335 16635 38341
rect 16577 38301 16589 38335
rect 16623 38301 16635 38335
rect 16577 38295 16635 38301
rect 16669 38335 16727 38341
rect 16669 38301 16681 38335
rect 16715 38332 16727 38335
rect 16942 38332 16948 38344
rect 16715 38304 16948 38332
rect 16715 38301 16727 38304
rect 16669 38295 16727 38301
rect 16942 38292 16948 38304
rect 17000 38292 17006 38344
rect 17034 38292 17040 38344
rect 17092 38332 17098 38344
rect 17402 38332 17408 38344
rect 17092 38304 17408 38332
rect 17092 38292 17098 38304
rect 17402 38292 17408 38304
rect 17460 38332 17466 38344
rect 17696 38341 17724 38372
rect 17788 38372 18236 38400
rect 17788 38341 17816 38372
rect 18230 38360 18236 38372
rect 18288 38360 18294 38412
rect 18340 38400 18368 38440
rect 19426 38428 19432 38480
rect 19484 38468 19490 38480
rect 19981 38471 20039 38477
rect 19981 38468 19993 38471
rect 19484 38440 19993 38468
rect 19484 38428 19490 38440
rect 19981 38437 19993 38440
rect 20027 38437 20039 38471
rect 19981 38431 20039 38437
rect 20993 38471 21051 38477
rect 20993 38437 21005 38471
rect 21039 38468 21051 38471
rect 22186 38468 22192 38480
rect 21039 38440 22192 38468
rect 21039 38437 21051 38440
rect 20993 38431 21051 38437
rect 22186 38428 22192 38440
rect 22244 38428 22250 38480
rect 22462 38468 22468 38480
rect 22388 38440 22468 38468
rect 22002 38400 22008 38412
rect 18340 38372 22008 38400
rect 22002 38360 22008 38372
rect 22060 38360 22066 38412
rect 17589 38335 17647 38341
rect 17589 38332 17601 38335
rect 17460 38304 17601 38332
rect 17460 38292 17466 38304
rect 17589 38301 17601 38304
rect 17635 38301 17647 38335
rect 17589 38295 17647 38301
rect 17681 38335 17739 38341
rect 17681 38301 17693 38335
rect 17727 38301 17739 38335
rect 17681 38295 17739 38301
rect 17773 38335 17831 38341
rect 17773 38301 17785 38335
rect 17819 38301 17831 38335
rect 17773 38295 17831 38301
rect 17957 38335 18015 38341
rect 17957 38301 17969 38335
rect 18003 38332 18015 38335
rect 18046 38332 18052 38344
rect 18003 38304 18052 38332
rect 18003 38301 18015 38304
rect 17957 38295 18015 38301
rect 12710 38224 12716 38276
rect 12768 38264 12774 38276
rect 13081 38267 13139 38273
rect 13081 38264 13093 38267
rect 12768 38236 13093 38264
rect 12768 38224 12774 38236
rect 13081 38233 13093 38236
rect 13127 38264 13139 38267
rect 14642 38264 14648 38276
rect 13127 38236 14648 38264
rect 13127 38233 13139 38236
rect 13081 38227 13139 38233
rect 14642 38224 14648 38236
rect 14700 38224 14706 38276
rect 15473 38267 15531 38273
rect 15473 38233 15485 38267
rect 15519 38233 15531 38267
rect 16482 38264 16488 38276
rect 16443 38236 16488 38264
rect 15473 38227 15531 38233
rect 11790 38156 11796 38208
rect 11848 38196 11854 38208
rect 12526 38196 12532 38208
rect 11848 38168 12532 38196
rect 11848 38156 11854 38168
rect 12526 38156 12532 38168
rect 12584 38196 12590 38208
rect 13281 38199 13339 38205
rect 13281 38196 13293 38199
rect 12584 38168 13293 38196
rect 12584 38156 12590 38168
rect 13281 38165 13293 38168
rect 13327 38165 13339 38199
rect 13446 38196 13452 38208
rect 13407 38168 13452 38196
rect 13281 38159 13339 38165
rect 13446 38156 13452 38168
rect 13504 38156 13510 38208
rect 14093 38199 14151 38205
rect 14093 38165 14105 38199
rect 14139 38196 14151 38199
rect 14366 38196 14372 38208
rect 14139 38168 14372 38196
rect 14139 38165 14151 38168
rect 14093 38159 14151 38165
rect 14366 38156 14372 38168
rect 14424 38156 14430 38208
rect 15488 38196 15516 38227
rect 16482 38224 16488 38236
rect 16540 38224 16546 38276
rect 16758 38264 16764 38276
rect 16592 38236 16764 38264
rect 16592 38196 16620 38236
rect 16758 38224 16764 38236
rect 16816 38224 16822 38276
rect 16850 38196 16856 38208
rect 15488 38168 16620 38196
rect 16811 38168 16856 38196
rect 16850 38156 16856 38168
rect 16908 38156 16914 38208
rect 17696 38196 17724 38295
rect 18046 38292 18052 38304
rect 18104 38332 18110 38344
rect 18874 38332 18880 38344
rect 18104 38304 18880 38332
rect 18104 38292 18110 38304
rect 18874 38292 18880 38304
rect 18932 38292 18938 38344
rect 19334 38292 19340 38344
rect 19392 38332 19398 38344
rect 19429 38335 19487 38341
rect 19429 38332 19441 38335
rect 19392 38304 19441 38332
rect 19392 38292 19398 38304
rect 19429 38301 19441 38304
rect 19475 38301 19487 38335
rect 19429 38295 19487 38301
rect 19536 38304 20208 38332
rect 17862 38224 17868 38276
rect 17920 38264 17926 38276
rect 19536 38264 19564 38304
rect 17920 38236 19564 38264
rect 19797 38267 19855 38273
rect 17920 38224 17926 38236
rect 19797 38233 19809 38267
rect 19843 38264 19855 38267
rect 20070 38264 20076 38276
rect 19843 38236 20076 38264
rect 19843 38233 19855 38236
rect 19797 38227 19855 38233
rect 20070 38224 20076 38236
rect 20128 38224 20134 38276
rect 20180 38264 20208 38304
rect 20714 38292 20720 38344
rect 20772 38332 20778 38344
rect 21266 38332 21272 38344
rect 20772 38304 21272 38332
rect 20772 38292 20778 38304
rect 21266 38292 21272 38304
rect 21324 38292 21330 38344
rect 21361 38335 21419 38341
rect 21361 38301 21373 38335
rect 21407 38301 21419 38335
rect 21361 38295 21419 38301
rect 20990 38264 20996 38276
rect 20180 38236 20996 38264
rect 20990 38224 20996 38236
rect 21048 38224 21054 38276
rect 21376 38264 21404 38295
rect 21450 38292 21456 38344
rect 21508 38332 21514 38344
rect 21637 38335 21695 38341
rect 21508 38304 21553 38332
rect 21508 38292 21514 38304
rect 21637 38301 21649 38335
rect 21683 38332 21695 38335
rect 21818 38332 21824 38344
rect 21683 38304 21824 38332
rect 21683 38301 21695 38304
rect 21637 38295 21695 38301
rect 21818 38292 21824 38304
rect 21876 38292 21882 38344
rect 21910 38292 21916 38344
rect 21968 38332 21974 38344
rect 22388 38341 22416 38440
rect 22462 38428 22468 38440
rect 22520 38428 22526 38480
rect 25130 38468 25136 38480
rect 25091 38440 25136 38468
rect 25130 38428 25136 38440
rect 25188 38428 25194 38480
rect 25685 38471 25743 38477
rect 25685 38437 25697 38471
rect 25731 38468 25743 38471
rect 26418 38468 26424 38480
rect 25731 38440 26424 38468
rect 25731 38437 25743 38440
rect 25685 38431 25743 38437
rect 26418 38428 26424 38440
rect 26476 38428 26482 38480
rect 22373 38335 22431 38341
rect 22373 38332 22385 38335
rect 21968 38304 22385 38332
rect 21968 38292 21974 38304
rect 22373 38301 22385 38304
rect 22419 38301 22431 38335
rect 22465 38335 22523 38341
rect 22465 38329 22477 38335
rect 22373 38295 22431 38301
rect 22460 38301 22477 38329
rect 22511 38301 22523 38335
rect 22460 38295 22523 38301
rect 22460 38264 22488 38295
rect 22554 38292 22560 38344
rect 22612 38332 22618 38344
rect 22741 38335 22799 38341
rect 22612 38304 22657 38332
rect 22612 38292 22618 38304
rect 22741 38301 22753 38335
rect 22787 38332 22799 38335
rect 23106 38332 23112 38344
rect 22787 38304 23112 38332
rect 22787 38301 22799 38304
rect 22741 38295 22799 38301
rect 23106 38292 23112 38304
rect 23164 38292 23170 38344
rect 23201 38335 23259 38341
rect 23201 38301 23213 38335
rect 23247 38301 23259 38335
rect 23201 38295 23259 38301
rect 23385 38335 23443 38341
rect 23385 38301 23397 38335
rect 23431 38332 23443 38335
rect 23750 38332 23756 38344
rect 23431 38304 23756 38332
rect 23431 38301 23443 38304
rect 23385 38295 23443 38301
rect 21100 38236 22488 38264
rect 21100 38208 21128 38236
rect 22830 38224 22836 38276
rect 22888 38264 22894 38276
rect 23216 38264 23244 38295
rect 22888 38236 23244 38264
rect 22888 38224 22894 38236
rect 21082 38196 21088 38208
rect 17696 38168 21088 38196
rect 21082 38156 21088 38168
rect 21140 38156 21146 38208
rect 22002 38156 22008 38208
rect 22060 38196 22066 38208
rect 23400 38196 23428 38295
rect 23750 38292 23756 38304
rect 23808 38292 23814 38344
rect 26050 38292 26056 38344
rect 26108 38332 26114 38344
rect 26145 38335 26203 38341
rect 26145 38332 26157 38335
rect 26108 38304 26157 38332
rect 26108 38292 26114 38304
rect 26145 38301 26157 38304
rect 26191 38301 26203 38335
rect 26326 38332 26332 38344
rect 26287 38304 26332 38332
rect 26145 38295 26203 38301
rect 26326 38292 26332 38304
rect 26384 38292 26390 38344
rect 25501 38267 25559 38273
rect 25501 38233 25513 38267
rect 25547 38264 25559 38267
rect 26237 38267 26295 38273
rect 26237 38264 26249 38267
rect 25547 38236 26249 38264
rect 25547 38233 25559 38236
rect 25501 38227 25559 38233
rect 26237 38233 26249 38236
rect 26283 38233 26295 38267
rect 26237 38227 26295 38233
rect 22060 38168 23428 38196
rect 22060 38156 22066 38168
rect 1104 38106 38824 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 38824 38106
rect 1104 38032 38824 38054
rect 10686 37992 10692 38004
rect 10647 37964 10692 37992
rect 10686 37952 10692 37964
rect 10744 37952 10750 38004
rect 12342 37952 12348 38004
rect 12400 37992 12406 38004
rect 12897 37995 12955 38001
rect 12897 37992 12909 37995
rect 12400 37964 12909 37992
rect 12400 37952 12406 37964
rect 12897 37961 12909 37964
rect 12943 37961 12955 37995
rect 14274 37992 14280 38004
rect 14235 37964 14280 37992
rect 12897 37955 12955 37961
rect 14274 37952 14280 37964
rect 14332 37952 14338 38004
rect 16206 37952 16212 38004
rect 16264 37992 16270 38004
rect 16482 37992 16488 38004
rect 16264 37964 16488 37992
rect 16264 37952 16270 37964
rect 16482 37952 16488 37964
rect 16540 37992 16546 38004
rect 18414 37992 18420 38004
rect 16540 37964 18420 37992
rect 16540 37952 16546 37964
rect 18414 37952 18420 37964
rect 18472 37952 18478 38004
rect 19334 37952 19340 38004
rect 19392 37992 19398 38004
rect 19429 37995 19487 38001
rect 19429 37992 19441 37995
rect 19392 37964 19441 37992
rect 19392 37952 19398 37964
rect 19429 37961 19441 37964
rect 19475 37961 19487 37995
rect 20070 37992 20076 38004
rect 20031 37964 20076 37992
rect 19429 37955 19487 37961
rect 20070 37952 20076 37964
rect 20128 37952 20134 38004
rect 21082 37952 21088 38004
rect 21140 37992 21146 38004
rect 21177 37995 21235 38001
rect 21177 37992 21189 37995
rect 21140 37964 21189 37992
rect 21140 37952 21146 37964
rect 21177 37961 21189 37964
rect 21223 37961 21235 37995
rect 21177 37955 21235 37961
rect 22189 37995 22247 38001
rect 22189 37961 22201 37995
rect 22235 37992 22247 37995
rect 22554 37992 22560 38004
rect 22235 37964 22560 37992
rect 22235 37961 22247 37964
rect 22189 37955 22247 37961
rect 22554 37952 22560 37964
rect 22612 37952 22618 38004
rect 25130 37952 25136 38004
rect 25188 37992 25194 38004
rect 25225 37995 25283 38001
rect 25225 37992 25237 37995
rect 25188 37964 25237 37992
rect 25188 37952 25194 37964
rect 25225 37961 25237 37964
rect 25271 37961 25283 37995
rect 27706 37992 27712 38004
rect 27667 37964 27712 37992
rect 25225 37955 25283 37961
rect 27706 37952 27712 37964
rect 27764 37952 27770 38004
rect 28350 37952 28356 38004
rect 28408 37992 28414 38004
rect 29381 37995 29439 38001
rect 29381 37992 29393 37995
rect 28408 37964 29393 37992
rect 28408 37952 28414 37964
rect 29381 37961 29393 37964
rect 29427 37961 29439 37995
rect 29381 37955 29439 37961
rect 12434 37924 12440 37936
rect 9324 37896 12440 37924
rect 8938 37816 8944 37868
rect 8996 37856 9002 37868
rect 9324 37865 9352 37896
rect 9582 37865 9588 37868
rect 9309 37859 9367 37865
rect 9309 37856 9321 37859
rect 8996 37828 9321 37856
rect 8996 37816 9002 37828
rect 9309 37825 9321 37828
rect 9355 37825 9367 37859
rect 9309 37819 9367 37825
rect 9576 37819 9588 37865
rect 9640 37856 9646 37868
rect 11532 37865 11560 37896
rect 12434 37884 12440 37896
rect 12492 37884 12498 37936
rect 14090 37924 14096 37936
rect 14051 37896 14096 37924
rect 14090 37884 14096 37896
rect 14148 37884 14154 37936
rect 14642 37884 14648 37936
rect 14700 37924 14706 37936
rect 14737 37927 14795 37933
rect 14737 37924 14749 37927
rect 14700 37896 14749 37924
rect 14700 37884 14706 37896
rect 14737 37893 14749 37896
rect 14783 37893 14795 37927
rect 14937 37927 14995 37933
rect 14937 37924 14949 37927
rect 14737 37887 14795 37893
rect 14844 37896 14949 37924
rect 11517 37859 11575 37865
rect 9640 37828 9676 37856
rect 9582 37816 9588 37819
rect 9640 37816 9646 37828
rect 11517 37825 11529 37859
rect 11563 37825 11575 37859
rect 11517 37819 11575 37825
rect 11606 37816 11612 37868
rect 11664 37856 11670 37868
rect 11773 37859 11831 37865
rect 11773 37856 11785 37859
rect 11664 37828 11785 37856
rect 11664 37816 11670 37828
rect 11773 37825 11785 37828
rect 11819 37825 11831 37859
rect 11773 37819 11831 37825
rect 13630 37816 13636 37868
rect 13688 37856 13694 37868
rect 14844 37856 14872 37896
rect 14937 37893 14949 37896
rect 14983 37893 14995 37927
rect 18506 37924 18512 37936
rect 18467 37896 18512 37924
rect 14937 37887 14995 37893
rect 18506 37884 18512 37896
rect 18564 37884 18570 37936
rect 19536 37896 20208 37924
rect 13688 37828 14872 37856
rect 16669 37859 16727 37865
rect 13688 37816 13694 37828
rect 16669 37825 16681 37859
rect 16715 37856 16727 37859
rect 18233 37859 18291 37865
rect 16715 37828 18184 37856
rect 16715 37825 16727 37828
rect 16669 37819 16727 37825
rect 16758 37748 16764 37800
rect 16816 37788 16822 37800
rect 16945 37791 17003 37797
rect 16945 37788 16957 37791
rect 16816 37760 16957 37788
rect 16816 37748 16822 37760
rect 16945 37757 16957 37760
rect 16991 37788 17003 37791
rect 17862 37788 17868 37800
rect 16991 37760 17868 37788
rect 16991 37757 17003 37760
rect 16945 37751 17003 37757
rect 17862 37748 17868 37760
rect 17920 37748 17926 37800
rect 18156 37788 18184 37828
rect 18233 37825 18245 37859
rect 18279 37856 18291 37859
rect 18322 37856 18328 37868
rect 18279 37828 18328 37856
rect 18279 37825 18291 37828
rect 18233 37819 18291 37825
rect 18322 37816 18328 37828
rect 18380 37816 18386 37868
rect 18414 37816 18420 37868
rect 18472 37856 18478 37868
rect 18472 37828 18517 37856
rect 18472 37816 18478 37828
rect 18598 37816 18604 37868
rect 18656 37856 18662 37868
rect 19536 37865 19564 37896
rect 20180 37865 20208 37896
rect 20990 37884 20996 37936
rect 21048 37924 21054 37936
rect 21821 37927 21879 37933
rect 21821 37924 21833 37927
rect 21048 37896 21833 37924
rect 21048 37884 21054 37896
rect 21821 37893 21833 37896
rect 21867 37893 21879 37927
rect 21821 37887 21879 37893
rect 22094 37884 22100 37936
rect 22152 37924 22158 37936
rect 22830 37924 22836 37936
rect 22152 37896 22836 37924
rect 22152 37884 22158 37896
rect 22830 37884 22836 37896
rect 22888 37884 22894 37936
rect 27890 37884 27896 37936
rect 27948 37924 27954 37936
rect 29181 37927 29239 37933
rect 29181 37924 29193 37927
rect 27948 37896 29193 37924
rect 27948 37884 27954 37896
rect 29181 37893 29193 37896
rect 29227 37893 29239 37927
rect 29181 37887 29239 37893
rect 19337 37859 19395 37865
rect 18656 37828 18701 37856
rect 18656 37816 18662 37828
rect 19337 37825 19349 37859
rect 19383 37825 19395 37859
rect 19337 37819 19395 37825
rect 19521 37859 19579 37865
rect 19521 37825 19533 37859
rect 19567 37825 19579 37859
rect 19521 37819 19579 37825
rect 19981 37859 20039 37865
rect 19981 37825 19993 37859
rect 20027 37825 20039 37859
rect 19981 37819 20039 37825
rect 20165 37859 20223 37865
rect 20165 37825 20177 37859
rect 20211 37856 20223 37859
rect 20622 37856 20628 37868
rect 20211 37828 20628 37856
rect 20211 37825 20223 37828
rect 20165 37819 20223 37825
rect 18506 37788 18512 37800
rect 18156 37760 18512 37788
rect 18506 37748 18512 37760
rect 18564 37748 18570 37800
rect 19352 37788 19380 37819
rect 19426 37788 19432 37800
rect 19339 37760 19432 37788
rect 19426 37748 19432 37760
rect 19484 37788 19490 37800
rect 19996 37788 20024 37819
rect 20622 37816 20628 37828
rect 20680 37816 20686 37868
rect 20806 37816 20812 37868
rect 20864 37856 20870 37868
rect 21085 37859 21143 37865
rect 21085 37856 21097 37859
rect 20864 37828 21097 37856
rect 20864 37816 20870 37828
rect 21085 37825 21097 37828
rect 21131 37825 21143 37859
rect 22002 37856 22008 37868
rect 21963 37828 22008 37856
rect 21085 37819 21143 37825
rect 22002 37816 22008 37828
rect 22060 37816 22066 37868
rect 25133 37859 25191 37865
rect 25133 37825 25145 37859
rect 25179 37825 25191 37859
rect 25133 37819 25191 37825
rect 19484 37760 20024 37788
rect 25148 37788 25176 37819
rect 25222 37816 25228 37868
rect 25280 37856 25286 37868
rect 25317 37859 25375 37865
rect 25317 37856 25329 37859
rect 25280 37828 25329 37856
rect 25280 37816 25286 37828
rect 25317 37825 25329 37828
rect 25363 37856 25375 37859
rect 26326 37856 26332 37868
rect 25363 37828 26332 37856
rect 25363 37825 25375 37828
rect 25317 37819 25375 37825
rect 26326 37816 26332 37828
rect 26384 37816 26390 37868
rect 27617 37859 27675 37865
rect 27617 37825 27629 37859
rect 27663 37856 27675 37859
rect 27663 37828 28764 37856
rect 27663 37825 27675 37828
rect 27617 37819 27675 37825
rect 26050 37788 26056 37800
rect 25148 37760 26056 37788
rect 19484 37748 19490 37760
rect 26050 37748 26056 37760
rect 26108 37748 26114 37800
rect 28261 37791 28319 37797
rect 28261 37757 28273 37791
rect 28307 37788 28319 37791
rect 28350 37788 28356 37800
rect 28307 37760 28356 37788
rect 28307 37757 28319 37760
rect 28261 37751 28319 37757
rect 28350 37748 28356 37760
rect 28408 37748 28414 37800
rect 28736 37797 28764 37828
rect 28721 37791 28779 37797
rect 28721 37757 28733 37791
rect 28767 37757 28779 37791
rect 28721 37751 28779 37757
rect 13722 37720 13728 37732
rect 13683 37692 13728 37720
rect 13722 37680 13728 37692
rect 13780 37680 13786 37732
rect 15105 37723 15163 37729
rect 15105 37720 15117 37723
rect 14108 37692 15117 37720
rect 14108 37661 14136 37692
rect 15105 37689 15117 37692
rect 15151 37689 15163 37723
rect 28166 37720 28172 37732
rect 15105 37683 15163 37689
rect 18156 37692 28172 37720
rect 14093 37655 14151 37661
rect 14093 37621 14105 37655
rect 14139 37621 14151 37655
rect 14093 37615 14151 37621
rect 14921 37655 14979 37661
rect 14921 37621 14933 37655
rect 14967 37652 14979 37655
rect 18156 37652 18184 37692
rect 28166 37680 28172 37692
rect 28224 37680 28230 37732
rect 28534 37720 28540 37732
rect 28495 37692 28540 37720
rect 28534 37680 28540 37692
rect 28592 37680 28598 37732
rect 37458 37720 37464 37732
rect 29380 37692 37464 37720
rect 14967 37624 18184 37652
rect 14967 37621 14979 37624
rect 14921 37615 14979 37621
rect 18230 37612 18236 37664
rect 18288 37652 18294 37664
rect 18785 37655 18843 37661
rect 18785 37652 18797 37655
rect 18288 37624 18797 37652
rect 18288 37612 18294 37624
rect 18785 37621 18797 37624
rect 18831 37621 18843 37655
rect 18785 37615 18843 37621
rect 18874 37612 18880 37664
rect 18932 37652 18938 37664
rect 21818 37652 21824 37664
rect 18932 37624 21824 37652
rect 18932 37612 18938 37624
rect 21818 37612 21824 37624
rect 21876 37612 21882 37664
rect 29380 37661 29408 37692
rect 37458 37680 37464 37692
rect 37516 37680 37522 37732
rect 29365 37655 29423 37661
rect 29365 37621 29377 37655
rect 29411 37621 29423 37655
rect 29546 37652 29552 37664
rect 29507 37624 29552 37652
rect 29365 37615 29423 37621
rect 29546 37612 29552 37624
rect 29604 37612 29610 37664
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 12069 37451 12127 37457
rect 12069 37417 12081 37451
rect 12115 37448 12127 37451
rect 13446 37448 13452 37460
rect 12115 37420 13452 37448
rect 12115 37417 12127 37420
rect 12069 37411 12127 37417
rect 13446 37408 13452 37420
rect 13504 37408 13510 37460
rect 16132 37420 16896 37448
rect 11701 37383 11759 37389
rect 11701 37349 11713 37383
rect 11747 37380 11759 37383
rect 11882 37380 11888 37392
rect 11747 37352 11888 37380
rect 11747 37349 11759 37352
rect 11701 37343 11759 37349
rect 11882 37340 11888 37352
rect 11940 37340 11946 37392
rect 13357 37383 13415 37389
rect 13357 37349 13369 37383
rect 13403 37380 13415 37383
rect 13722 37380 13728 37392
rect 13403 37352 13728 37380
rect 13403 37349 13415 37352
rect 13357 37343 13415 37349
rect 13722 37340 13728 37352
rect 13780 37340 13786 37392
rect 15654 37340 15660 37392
rect 15712 37380 15718 37392
rect 16132 37380 16160 37420
rect 16574 37380 16580 37392
rect 15712 37352 16160 37380
rect 15712 37340 15718 37352
rect 8938 37312 8944 37324
rect 8899 37284 8944 37312
rect 8938 37272 8944 37284
rect 8996 37272 9002 37324
rect 16022 37312 16028 37324
rect 15983 37284 16028 37312
rect 16022 37272 16028 37284
rect 16080 37272 16086 37324
rect 13262 37204 13268 37256
rect 13320 37244 13326 37256
rect 14093 37247 14151 37253
rect 14093 37244 14105 37247
rect 13320 37216 14105 37244
rect 13320 37204 13326 37216
rect 14093 37213 14105 37216
rect 14139 37244 14151 37247
rect 15746 37244 15752 37256
rect 14139 37216 15752 37244
rect 14139 37213 14151 37216
rect 14093 37207 14151 37213
rect 15746 37204 15752 37216
rect 15804 37204 15810 37256
rect 16132 37244 16160 37352
rect 16408 37352 16580 37380
rect 16209 37247 16267 37253
rect 16209 37244 16221 37247
rect 16132 37216 16221 37244
rect 16209 37213 16221 37216
rect 16255 37213 16267 37247
rect 16209 37207 16267 37213
rect 16301 37247 16359 37253
rect 16301 37213 16313 37247
rect 16347 37244 16359 37247
rect 16408 37244 16436 37352
rect 16574 37340 16580 37352
rect 16632 37340 16638 37392
rect 16868 37312 16896 37420
rect 16942 37408 16948 37460
rect 17000 37448 17006 37460
rect 18598 37448 18604 37460
rect 17000 37420 18604 37448
rect 17000 37408 17006 37420
rect 18598 37408 18604 37420
rect 18656 37408 18662 37460
rect 23661 37451 23719 37457
rect 23661 37417 23673 37451
rect 23707 37448 23719 37451
rect 24302 37448 24308 37460
rect 23707 37420 24308 37448
rect 23707 37417 23719 37420
rect 23661 37411 23719 37417
rect 24302 37408 24308 37420
rect 24360 37408 24366 37460
rect 23290 37380 23296 37392
rect 23251 37352 23296 37380
rect 23290 37340 23296 37352
rect 23348 37340 23354 37392
rect 23382 37340 23388 37392
rect 23440 37380 23446 37392
rect 24949 37383 25007 37389
rect 24949 37380 24961 37383
rect 23440 37352 24961 37380
rect 23440 37340 23446 37352
rect 24949 37349 24961 37352
rect 24995 37349 25007 37383
rect 24949 37343 25007 37349
rect 17678 37312 17684 37324
rect 16868 37284 16988 37312
rect 17639 37284 17684 37312
rect 16347 37216 16436 37244
rect 16485 37247 16543 37253
rect 16347 37213 16359 37216
rect 16301 37207 16359 37213
rect 16485 37213 16497 37247
rect 16531 37213 16543 37247
rect 16485 37207 16543 37213
rect 16572 37247 16630 37253
rect 16572 37213 16584 37247
rect 16618 37244 16630 37247
rect 16850 37244 16856 37256
rect 16618 37216 16856 37244
rect 16618 37213 16630 37216
rect 16572 37207 16630 37213
rect 9208 37179 9266 37185
rect 9208 37145 9220 37179
rect 9254 37176 9266 37179
rect 9398 37176 9404 37188
rect 9254 37148 9404 37176
rect 9254 37145 9266 37148
rect 9208 37139 9266 37145
rect 9398 37136 9404 37148
rect 9456 37136 9462 37188
rect 12989 37179 13047 37185
rect 12989 37145 13001 37179
rect 13035 37176 13047 37179
rect 13630 37176 13636 37188
rect 13035 37148 13636 37176
rect 13035 37145 13047 37148
rect 12989 37139 13047 37145
rect 13630 37136 13636 37148
rect 13688 37136 13694 37188
rect 14366 37185 14372 37188
rect 14360 37176 14372 37185
rect 14327 37148 14372 37176
rect 14360 37139 14372 37148
rect 14366 37136 14372 37139
rect 14424 37136 14430 37188
rect 14642 37136 14648 37188
rect 14700 37176 14706 37188
rect 16500 37176 16528 37207
rect 16850 37204 16856 37216
rect 16908 37204 16914 37256
rect 16960 37244 16988 37284
rect 17678 37272 17684 37284
rect 17736 37272 17742 37324
rect 28902 37312 28908 37324
rect 19306 37284 21128 37312
rect 17865 37247 17923 37253
rect 17865 37244 17877 37247
rect 16960 37216 17877 37244
rect 17865 37213 17877 37216
rect 17911 37213 17923 37247
rect 17865 37207 17923 37213
rect 16666 37176 16672 37188
rect 14700 37148 15700 37176
rect 16500 37148 16672 37176
rect 14700 37136 14706 37148
rect 10318 37108 10324 37120
rect 10279 37080 10324 37108
rect 10318 37068 10324 37080
rect 10376 37068 10382 37120
rect 11882 37068 11888 37120
rect 11940 37108 11946 37120
rect 12069 37111 12127 37117
rect 12069 37108 12081 37111
rect 11940 37080 12081 37108
rect 11940 37068 11946 37080
rect 12069 37077 12081 37080
rect 12115 37077 12127 37111
rect 12250 37108 12256 37120
rect 12211 37080 12256 37108
rect 12069 37071 12127 37077
rect 12250 37068 12256 37080
rect 12308 37068 12314 37120
rect 13449 37111 13507 37117
rect 13449 37077 13461 37111
rect 13495 37108 13507 37111
rect 13538 37108 13544 37120
rect 13495 37080 13544 37108
rect 13495 37077 13507 37080
rect 13449 37071 13507 37077
rect 13538 37068 13544 37080
rect 13596 37068 13602 37120
rect 15473 37111 15531 37117
rect 15473 37077 15485 37111
rect 15519 37108 15531 37111
rect 15562 37108 15568 37120
rect 15519 37080 15568 37108
rect 15519 37077 15531 37080
rect 15473 37071 15531 37077
rect 15562 37068 15568 37080
rect 15620 37068 15626 37120
rect 15672 37108 15700 37148
rect 16666 37136 16672 37148
rect 16724 37136 16730 37188
rect 17880 37176 17908 37207
rect 17954 37204 17960 37256
rect 18012 37244 18018 37256
rect 18138 37244 18144 37256
rect 18012 37216 18057 37244
rect 18099 37216 18144 37244
rect 18012 37204 18018 37216
rect 18138 37204 18144 37216
rect 18196 37204 18202 37256
rect 18230 37204 18236 37256
rect 18288 37244 18294 37256
rect 18288 37216 18333 37244
rect 18288 37204 18294 37216
rect 18598 37204 18604 37256
rect 18656 37244 18662 37256
rect 19306 37244 19334 37284
rect 18656 37216 19334 37244
rect 20901 37247 20959 37253
rect 18656 37204 18662 37216
rect 20901 37213 20913 37247
rect 20947 37244 20959 37247
rect 20990 37244 20996 37256
rect 20947 37216 20996 37244
rect 20947 37213 20959 37216
rect 20901 37207 20959 37213
rect 20990 37204 20996 37216
rect 21048 37204 21054 37256
rect 21100 37244 21128 37284
rect 26436 37284 28908 37312
rect 21269 37247 21327 37253
rect 21269 37244 21281 37247
rect 21100 37216 21281 37244
rect 21269 37213 21281 37216
rect 21315 37244 21327 37247
rect 22186 37244 22192 37256
rect 21315 37216 22192 37244
rect 21315 37213 21327 37216
rect 21269 37207 21327 37213
rect 22186 37204 22192 37216
rect 22244 37204 22250 37256
rect 25038 37204 25044 37256
rect 25096 37244 25102 37256
rect 25409 37247 25467 37253
rect 25409 37244 25421 37247
rect 25096 37216 25421 37244
rect 25096 37204 25102 37216
rect 25409 37213 25421 37216
rect 25455 37244 25467 37247
rect 26436 37244 26464 37284
rect 28902 37272 28908 37284
rect 28960 37272 28966 37324
rect 27246 37244 27252 37256
rect 25455 37216 26464 37244
rect 27207 37216 27252 37244
rect 25455 37213 25467 37216
rect 25409 37207 25467 37213
rect 27246 37204 27252 37216
rect 27304 37204 27310 37256
rect 18322 37176 18328 37188
rect 17880 37148 18328 37176
rect 18322 37136 18328 37148
rect 18380 37136 18386 37188
rect 18414 37136 18420 37188
rect 18472 37176 18478 37188
rect 21082 37176 21088 37188
rect 18472 37148 21088 37176
rect 18472 37136 18478 37148
rect 21082 37136 21088 37148
rect 21140 37136 21146 37188
rect 21177 37179 21235 37185
rect 21177 37145 21189 37179
rect 21223 37176 21235 37179
rect 22094 37176 22100 37188
rect 21223 37148 22100 37176
rect 21223 37145 21235 37148
rect 21177 37139 21235 37145
rect 22094 37136 22100 37148
rect 22152 37136 22158 37188
rect 24765 37179 24823 37185
rect 24765 37145 24777 37179
rect 24811 37176 24823 37179
rect 25314 37176 25320 37188
rect 24811 37148 25320 37176
rect 24811 37145 24823 37148
rect 24765 37139 24823 37145
rect 25314 37136 25320 37148
rect 25372 37136 25378 37188
rect 25676 37179 25734 37185
rect 25676 37145 25688 37179
rect 25722 37176 25734 37179
rect 27614 37176 27620 37188
rect 25722 37148 27620 37176
rect 25722 37145 25734 37148
rect 25676 37139 25734 37145
rect 27614 37136 27620 37148
rect 27672 37136 27678 37188
rect 19150 37108 19156 37120
rect 15672 37080 19156 37108
rect 19150 37068 19156 37080
rect 19208 37068 19214 37120
rect 19334 37068 19340 37120
rect 19392 37108 19398 37120
rect 20162 37108 20168 37120
rect 19392 37080 20168 37108
rect 19392 37068 19398 37080
rect 20162 37068 20168 37080
rect 20220 37068 20226 37120
rect 20714 37068 20720 37120
rect 20772 37108 20778 37120
rect 21453 37111 21511 37117
rect 21453 37108 21465 37111
rect 20772 37080 21465 37108
rect 20772 37068 20778 37080
rect 21453 37077 21465 37080
rect 21499 37077 21511 37111
rect 21453 37071 21511 37077
rect 23661 37111 23719 37117
rect 23661 37077 23673 37111
rect 23707 37108 23719 37111
rect 23750 37108 23756 37120
rect 23707 37080 23756 37108
rect 23707 37077 23719 37080
rect 23661 37071 23719 37077
rect 23750 37068 23756 37080
rect 23808 37068 23814 37120
rect 23845 37111 23903 37117
rect 23845 37077 23857 37111
rect 23891 37108 23903 37111
rect 24486 37108 24492 37120
rect 23891 37080 24492 37108
rect 23891 37077 23903 37080
rect 23845 37071 23903 37077
rect 24486 37068 24492 37080
rect 24544 37068 24550 37120
rect 26786 37108 26792 37120
rect 26747 37080 26792 37108
rect 26786 37068 26792 37080
rect 26844 37068 26850 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 11882 36904 11888 36916
rect 11843 36876 11888 36904
rect 11882 36864 11888 36876
rect 11940 36864 11946 36916
rect 13449 36907 13507 36913
rect 13449 36873 13461 36907
rect 13495 36904 13507 36907
rect 13722 36904 13728 36916
rect 13495 36876 13728 36904
rect 13495 36873 13507 36876
rect 13449 36867 13507 36873
rect 13722 36864 13728 36876
rect 13780 36864 13786 36916
rect 14090 36904 14096 36916
rect 14051 36876 14096 36904
rect 14090 36864 14096 36876
rect 14148 36864 14154 36916
rect 16666 36864 16672 36916
rect 16724 36904 16730 36916
rect 17037 36907 17095 36913
rect 17037 36904 17049 36907
rect 16724 36876 17049 36904
rect 16724 36864 16730 36876
rect 17037 36873 17049 36876
rect 17083 36873 17095 36907
rect 18690 36904 18696 36916
rect 18651 36876 18696 36904
rect 17037 36867 17095 36873
rect 18690 36864 18696 36876
rect 18748 36864 18754 36916
rect 22370 36904 22376 36916
rect 20456 36876 22376 36904
rect 15749 36839 15807 36845
rect 11900 36808 12572 36836
rect 8938 36728 8944 36780
rect 8996 36768 9002 36780
rect 9858 36777 9864 36780
rect 9585 36771 9643 36777
rect 9585 36768 9597 36771
rect 8996 36740 9597 36768
rect 8996 36728 9002 36740
rect 9585 36737 9597 36740
rect 9631 36737 9643 36771
rect 9585 36731 9643 36737
rect 9852 36731 9864 36777
rect 9916 36768 9922 36780
rect 11900 36777 11928 36808
rect 12544 36780 12572 36808
rect 13556 36808 14228 36836
rect 11701 36771 11759 36777
rect 9916 36740 9952 36768
rect 9858 36728 9864 36731
rect 9916 36728 9922 36740
rect 11701 36737 11713 36771
rect 11747 36737 11759 36771
rect 11701 36731 11759 36737
rect 11885 36771 11943 36777
rect 11885 36737 11897 36771
rect 11931 36737 11943 36771
rect 11885 36731 11943 36737
rect 12345 36771 12403 36777
rect 12345 36737 12357 36771
rect 12391 36768 12403 36771
rect 12526 36768 12532 36780
rect 12391 36740 12425 36768
rect 12487 36740 12532 36768
rect 12391 36737 12403 36740
rect 12345 36731 12403 36737
rect 11716 36700 11744 36731
rect 12360 36700 12388 36731
rect 12526 36728 12532 36740
rect 12584 36728 12590 36780
rect 13556 36777 13584 36808
rect 14200 36777 14228 36808
rect 15749 36805 15761 36839
rect 15795 36836 15807 36839
rect 16206 36836 16212 36848
rect 15795 36808 16212 36836
rect 15795 36805 15807 36808
rect 15749 36799 15807 36805
rect 16206 36796 16212 36808
rect 16264 36796 16270 36848
rect 16942 36836 16948 36848
rect 16776 36808 16948 36836
rect 13357 36771 13415 36777
rect 13357 36737 13369 36771
rect 13403 36737 13415 36771
rect 13357 36731 13415 36737
rect 13541 36771 13599 36777
rect 13541 36737 13553 36771
rect 13587 36737 13599 36771
rect 13541 36731 13599 36737
rect 14001 36771 14059 36777
rect 14001 36737 14013 36771
rect 14047 36737 14059 36771
rect 14001 36731 14059 36737
rect 14185 36771 14243 36777
rect 14185 36737 14197 36771
rect 14231 36737 14243 36771
rect 15562 36768 15568 36780
rect 15523 36740 15568 36768
rect 14185 36731 14243 36737
rect 12802 36700 12808 36712
rect 11716 36672 12808 36700
rect 12802 36660 12808 36672
rect 12860 36660 12866 36712
rect 13372 36700 13400 36731
rect 13814 36700 13820 36712
rect 13372 36672 13820 36700
rect 13814 36660 13820 36672
rect 13872 36700 13878 36712
rect 14016 36700 14044 36731
rect 13872 36672 14044 36700
rect 13872 36660 13878 36672
rect 11974 36592 11980 36644
rect 12032 36632 12038 36644
rect 12345 36635 12403 36641
rect 12345 36632 12357 36635
rect 12032 36604 12357 36632
rect 12032 36592 12038 36604
rect 12345 36601 12357 36604
rect 12391 36601 12403 36635
rect 14200 36632 14228 36731
rect 15562 36728 15568 36740
rect 15620 36728 15626 36780
rect 15841 36771 15899 36777
rect 15841 36737 15853 36771
rect 15887 36737 15899 36771
rect 15841 36731 15899 36737
rect 15933 36771 15991 36777
rect 15933 36737 15945 36771
rect 15979 36768 15991 36771
rect 16776 36768 16804 36808
rect 16942 36796 16948 36808
rect 17000 36796 17006 36848
rect 19150 36836 19156 36848
rect 19111 36808 19156 36836
rect 19150 36796 19156 36808
rect 19208 36796 19214 36848
rect 19353 36839 19411 36845
rect 19353 36836 19365 36839
rect 19260 36808 19365 36836
rect 15979 36740 16804 36768
rect 16853 36771 16911 36777
rect 15979 36737 15991 36740
rect 15933 36731 15991 36737
rect 16853 36737 16865 36771
rect 16899 36768 16911 36771
rect 17678 36768 17684 36780
rect 16899 36740 17684 36768
rect 16899 36737 16911 36740
rect 16853 36731 16911 36737
rect 15856 36700 15884 36731
rect 17678 36728 17684 36740
rect 17736 36728 17742 36780
rect 19260 36768 19288 36808
rect 19353 36805 19365 36808
rect 19399 36805 19411 36839
rect 19353 36799 19411 36805
rect 19886 36768 19892 36780
rect 18248 36740 19288 36768
rect 19352 36740 19892 36768
rect 16022 36700 16028 36712
rect 15856 36672 16028 36700
rect 16022 36660 16028 36672
rect 16080 36660 16086 36712
rect 16669 36703 16727 36709
rect 16669 36669 16681 36703
rect 16715 36700 16727 36703
rect 17586 36700 17592 36712
rect 16715 36672 17592 36700
rect 16715 36669 16727 36672
rect 16669 36663 16727 36669
rect 16684 36632 16712 36663
rect 17586 36660 17592 36672
rect 17644 36660 17650 36712
rect 17954 36660 17960 36712
rect 18012 36700 18018 36712
rect 18248 36709 18276 36740
rect 18233 36703 18291 36709
rect 18233 36700 18245 36703
rect 18012 36672 18245 36700
rect 18012 36660 18018 36672
rect 18233 36669 18245 36672
rect 18279 36669 18291 36703
rect 18233 36663 18291 36669
rect 18322 36660 18328 36712
rect 18380 36700 18386 36712
rect 19352 36700 19380 36740
rect 19886 36728 19892 36740
rect 19944 36768 19950 36780
rect 20456 36777 20484 36876
rect 22370 36864 22376 36876
rect 22428 36864 22434 36916
rect 23109 36907 23167 36913
rect 23109 36873 23121 36907
rect 23155 36904 23167 36907
rect 23290 36904 23296 36916
rect 23155 36876 23296 36904
rect 23155 36873 23167 36876
rect 23109 36867 23167 36873
rect 23290 36864 23296 36876
rect 23348 36864 23354 36916
rect 23750 36904 23756 36916
rect 23711 36876 23756 36904
rect 23750 36864 23756 36876
rect 23808 36864 23814 36916
rect 26418 36904 26424 36916
rect 26379 36876 26424 36904
rect 26418 36864 26424 36876
rect 26476 36864 26482 36916
rect 27614 36904 27620 36916
rect 27575 36876 27620 36904
rect 27614 36864 27620 36876
rect 27672 36864 27678 36916
rect 29822 36904 29828 36916
rect 27724 36876 29828 36904
rect 26786 36836 26792 36848
rect 21836 36808 26792 36836
rect 20349 36771 20407 36777
rect 20349 36768 20361 36771
rect 19944 36740 20361 36768
rect 19944 36728 19950 36740
rect 20349 36737 20361 36740
rect 20395 36737 20407 36771
rect 20349 36731 20407 36737
rect 20441 36771 20499 36777
rect 20441 36737 20453 36771
rect 20487 36737 20499 36771
rect 20441 36731 20499 36737
rect 20625 36771 20683 36777
rect 20625 36737 20637 36771
rect 20671 36737 20683 36771
rect 20625 36731 20683 36737
rect 18380 36672 19380 36700
rect 20640 36700 20668 36731
rect 20714 36728 20720 36780
rect 20772 36768 20778 36780
rect 21836 36777 21864 36808
rect 26786 36796 26792 36808
rect 26844 36796 26850 36848
rect 21821 36771 21879 36777
rect 20772 36740 20817 36768
rect 20772 36728 20778 36740
rect 21821 36737 21833 36771
rect 21867 36737 21879 36771
rect 21821 36731 21879 36737
rect 22005 36771 22063 36777
rect 22005 36737 22017 36771
rect 22051 36737 22063 36771
rect 22005 36731 22063 36737
rect 22097 36771 22155 36777
rect 22097 36737 22109 36771
rect 22143 36737 22155 36771
rect 22097 36731 22155 36737
rect 20990 36700 20996 36712
rect 20640 36672 20996 36700
rect 18380 36660 18386 36672
rect 20990 36660 20996 36672
rect 21048 36660 21054 36712
rect 21082 36660 21088 36712
rect 21140 36700 21146 36712
rect 22020 36700 22048 36731
rect 21140 36672 22048 36700
rect 22112 36700 22140 36731
rect 22186 36728 22192 36780
rect 22244 36768 22250 36780
rect 23017 36771 23075 36777
rect 22244 36740 22289 36768
rect 22244 36728 22250 36740
rect 23017 36737 23029 36771
rect 23063 36768 23075 36771
rect 23201 36771 23259 36777
rect 23063 36740 23152 36768
rect 23063 36737 23075 36740
rect 23017 36731 23075 36737
rect 23124 36700 23152 36740
rect 23201 36737 23213 36771
rect 23247 36768 23259 36771
rect 23382 36768 23388 36780
rect 23247 36740 23388 36768
rect 23247 36737 23259 36740
rect 23201 36731 23259 36737
rect 23382 36728 23388 36740
rect 23440 36728 23446 36780
rect 23658 36768 23664 36780
rect 23619 36740 23664 36768
rect 23658 36728 23664 36740
rect 23716 36728 23722 36780
rect 23845 36771 23903 36777
rect 23845 36737 23857 36771
rect 23891 36737 23903 36771
rect 24486 36768 24492 36780
rect 24447 36740 24492 36768
rect 23845 36731 23903 36737
rect 22112 36672 23152 36700
rect 23400 36700 23428 36728
rect 23860 36700 23888 36731
rect 24486 36728 24492 36740
rect 24544 36728 24550 36780
rect 25038 36768 25044 36780
rect 24999 36740 25044 36768
rect 25038 36728 25044 36740
rect 25096 36728 25102 36780
rect 25308 36771 25366 36777
rect 25308 36737 25320 36771
rect 25354 36768 25366 36771
rect 26326 36768 26332 36780
rect 25354 36740 26332 36768
rect 25354 36737 25366 36740
rect 25308 36731 25366 36737
rect 26326 36728 26332 36740
rect 26384 36728 26390 36780
rect 23400 36672 23888 36700
rect 21140 36660 21146 36672
rect 14200 36604 16712 36632
rect 18601 36635 18659 36641
rect 12345 36595 12403 36601
rect 18601 36601 18613 36635
rect 18647 36632 18659 36635
rect 19242 36632 19248 36644
rect 18647 36604 19248 36632
rect 18647 36601 18659 36604
rect 18601 36595 18659 36601
rect 19242 36592 19248 36604
rect 19300 36592 19306 36644
rect 23124 36632 23152 36672
rect 23658 36632 23664 36644
rect 19352 36604 23060 36632
rect 23124 36604 23664 36632
rect 10965 36567 11023 36573
rect 10965 36533 10977 36567
rect 11011 36564 11023 36567
rect 11146 36564 11152 36576
rect 11011 36536 11152 36564
rect 11011 36533 11023 36536
rect 10965 36527 11023 36533
rect 11146 36524 11152 36536
rect 11204 36564 11210 36576
rect 11698 36564 11704 36576
rect 11204 36536 11704 36564
rect 11204 36524 11210 36536
rect 11698 36524 11704 36536
rect 11756 36524 11762 36576
rect 15838 36524 15844 36576
rect 15896 36564 15902 36576
rect 19352 36573 19380 36604
rect 16117 36567 16175 36573
rect 16117 36564 16129 36567
rect 15896 36536 16129 36564
rect 15896 36524 15902 36536
rect 16117 36533 16129 36536
rect 16163 36533 16175 36567
rect 16117 36527 16175 36533
rect 19337 36567 19395 36573
rect 19337 36533 19349 36567
rect 19383 36533 19395 36567
rect 19337 36527 19395 36533
rect 19521 36567 19579 36573
rect 19521 36533 19533 36567
rect 19567 36564 19579 36567
rect 19610 36564 19616 36576
rect 19567 36536 19616 36564
rect 19567 36533 19579 36536
rect 19521 36527 19579 36533
rect 19610 36524 19616 36536
rect 19668 36524 19674 36576
rect 20162 36564 20168 36576
rect 20123 36536 20168 36564
rect 20162 36524 20168 36536
rect 20220 36524 20226 36576
rect 21358 36524 21364 36576
rect 21416 36564 21422 36576
rect 22373 36567 22431 36573
rect 22373 36564 22385 36567
rect 21416 36536 22385 36564
rect 21416 36524 21422 36536
rect 22373 36533 22385 36536
rect 22419 36533 22431 36567
rect 23032 36564 23060 36604
rect 23658 36592 23664 36604
rect 23716 36592 23722 36644
rect 23768 36604 25084 36632
rect 23768 36564 23796 36604
rect 24302 36564 24308 36576
rect 23032 36536 23796 36564
rect 24263 36536 24308 36564
rect 22373 36527 22431 36533
rect 24302 36524 24308 36536
rect 24360 36524 24366 36576
rect 25056 36564 25084 36604
rect 27724 36564 27752 36876
rect 29822 36864 29828 36876
rect 29880 36864 29886 36916
rect 28626 36836 28632 36848
rect 28587 36808 28632 36836
rect 28626 36796 28632 36808
rect 28684 36796 28690 36848
rect 27801 36771 27859 36777
rect 27801 36737 27813 36771
rect 27847 36768 27859 36771
rect 27847 36740 28856 36768
rect 27847 36737 27859 36740
rect 27801 36731 27859 36737
rect 28261 36703 28319 36709
rect 28261 36669 28273 36703
rect 28307 36700 28319 36703
rect 28534 36700 28540 36712
rect 28307 36672 28540 36700
rect 28307 36669 28319 36672
rect 28261 36663 28319 36669
rect 28534 36660 28540 36672
rect 28592 36660 28598 36712
rect 28828 36641 28856 36740
rect 28813 36635 28871 36641
rect 28813 36601 28825 36635
rect 28859 36601 28871 36635
rect 28813 36595 28871 36601
rect 25056 36536 27752 36564
rect 28629 36567 28687 36573
rect 28629 36533 28641 36567
rect 28675 36564 28687 36567
rect 29546 36564 29552 36576
rect 28675 36536 29552 36564
rect 28675 36533 28687 36536
rect 28629 36527 28687 36533
rect 29546 36524 29552 36536
rect 29604 36524 29610 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 13170 36360 13176 36372
rect 13131 36332 13176 36360
rect 13170 36320 13176 36332
rect 13228 36320 13234 36372
rect 16206 36360 16212 36372
rect 16167 36332 16212 36360
rect 16206 36320 16212 36332
rect 16264 36320 16270 36372
rect 16942 36360 16948 36372
rect 16903 36332 16948 36360
rect 16942 36320 16948 36332
rect 17000 36320 17006 36372
rect 18138 36320 18144 36372
rect 18196 36360 18202 36372
rect 18233 36363 18291 36369
rect 18233 36360 18245 36363
rect 18196 36332 18245 36360
rect 18196 36320 18202 36332
rect 18233 36329 18245 36332
rect 18279 36329 18291 36363
rect 19610 36360 19616 36372
rect 19571 36332 19616 36360
rect 18233 36323 18291 36329
rect 19610 36320 19616 36332
rect 19668 36320 19674 36372
rect 22281 36363 22339 36369
rect 22281 36329 22293 36363
rect 22327 36360 22339 36363
rect 25685 36363 25743 36369
rect 22327 36332 25636 36360
rect 22327 36329 22339 36332
rect 22281 36323 22339 36329
rect 19797 36295 19855 36301
rect 19797 36292 19809 36295
rect 12406 36264 19809 36292
rect 11793 36159 11851 36165
rect 11793 36125 11805 36159
rect 11839 36156 11851 36159
rect 12406 36156 12434 36264
rect 19797 36261 19809 36264
rect 19843 36261 19855 36295
rect 19797 36255 19855 36261
rect 19886 36252 19892 36304
rect 19944 36292 19950 36304
rect 22554 36292 22560 36304
rect 19944 36264 20852 36292
rect 19944 36252 19950 36264
rect 17865 36227 17923 36233
rect 17865 36193 17877 36227
rect 17911 36224 17923 36227
rect 18414 36224 18420 36236
rect 17911 36196 18420 36224
rect 17911 36193 17923 36196
rect 17865 36187 17923 36193
rect 18414 36184 18420 36196
rect 18472 36184 18478 36236
rect 19150 36184 19156 36236
rect 19208 36224 19214 36236
rect 19208 36196 20760 36224
rect 19208 36184 19214 36196
rect 11839 36128 12434 36156
rect 11839 36125 11851 36128
rect 11793 36119 11851 36125
rect 13078 36116 13084 36168
rect 13136 36156 13142 36168
rect 13173 36159 13231 36165
rect 13173 36156 13185 36159
rect 13136 36128 13185 36156
rect 13136 36116 13142 36128
rect 13173 36125 13185 36128
rect 13219 36125 13231 36159
rect 13173 36119 13231 36125
rect 13357 36159 13415 36165
rect 13357 36125 13369 36159
rect 13403 36156 13415 36159
rect 16022 36156 16028 36168
rect 13403 36128 16028 36156
rect 13403 36125 13415 36128
rect 13357 36119 13415 36125
rect 16022 36116 16028 36128
rect 16080 36116 16086 36168
rect 17678 36116 17684 36168
rect 17736 36156 17742 36168
rect 18049 36159 18107 36165
rect 18049 36156 18061 36159
rect 17736 36128 18061 36156
rect 17736 36116 17742 36128
rect 18049 36125 18061 36128
rect 18095 36125 18107 36159
rect 19242 36156 19248 36168
rect 19203 36128 19248 36156
rect 18049 36119 18107 36125
rect 19242 36116 19248 36128
rect 19300 36116 19306 36168
rect 15562 36048 15568 36100
rect 15620 36088 15626 36100
rect 16117 36091 16175 36097
rect 16117 36088 16129 36091
rect 15620 36060 16129 36088
rect 15620 36048 15626 36060
rect 16117 36057 16129 36060
rect 16163 36057 16175 36091
rect 16117 36051 16175 36057
rect 16853 36091 16911 36097
rect 16853 36057 16865 36091
rect 16899 36088 16911 36091
rect 17770 36088 17776 36100
rect 16899 36060 17776 36088
rect 16899 36057 16911 36060
rect 16853 36051 16911 36057
rect 17770 36048 17776 36060
rect 17828 36048 17834 36100
rect 19613 36091 19671 36097
rect 19613 36057 19625 36091
rect 19659 36088 19671 36091
rect 20622 36088 20628 36100
rect 19659 36060 20628 36088
rect 19659 36057 19671 36060
rect 19613 36051 19671 36057
rect 20622 36048 20628 36060
rect 20680 36048 20686 36100
rect 20732 36088 20760 36196
rect 20824 36156 20852 36264
rect 21100 36264 22560 36292
rect 21100 36165 21128 36264
rect 22554 36252 22560 36264
rect 22612 36252 22618 36304
rect 22094 36224 22100 36236
rect 21284 36196 22100 36224
rect 21284 36165 21312 36196
rect 22094 36184 22100 36196
rect 22152 36184 22158 36236
rect 25608 36224 25636 36332
rect 25685 36329 25697 36363
rect 25731 36360 25743 36363
rect 37274 36360 37280 36372
rect 25731 36332 37280 36360
rect 25731 36329 25743 36332
rect 25685 36323 25743 36329
rect 37274 36320 37280 36332
rect 37332 36320 37338 36372
rect 26326 36292 26332 36304
rect 26287 36264 26332 36292
rect 26326 36252 26332 36264
rect 26384 36252 26390 36304
rect 29914 36292 29920 36304
rect 28368 36264 29920 36292
rect 28368 36224 28396 36264
rect 29914 36252 29920 36264
rect 29972 36252 29978 36304
rect 28534 36224 28540 36236
rect 25608 36196 28396 36224
rect 28495 36196 28540 36224
rect 28534 36184 28540 36196
rect 28592 36184 28598 36236
rect 20993 36159 21051 36165
rect 20993 36156 21005 36159
rect 20824 36128 21005 36156
rect 20993 36125 21005 36128
rect 21039 36125 21051 36159
rect 20993 36119 21051 36125
rect 21085 36159 21143 36165
rect 21085 36125 21097 36159
rect 21131 36125 21143 36159
rect 21085 36119 21143 36125
rect 21269 36159 21327 36165
rect 21269 36125 21281 36159
rect 21315 36125 21327 36159
rect 21269 36119 21327 36125
rect 21358 36116 21364 36168
rect 21416 36156 21422 36168
rect 26510 36156 26516 36168
rect 21416 36128 21461 36156
rect 26471 36128 26516 36156
rect 21416 36116 21422 36128
rect 26510 36116 26516 36128
rect 26568 36116 26574 36168
rect 28442 36156 28448 36168
rect 28403 36128 28448 36156
rect 28442 36116 28448 36128
rect 28500 36116 28506 36168
rect 28629 36159 28687 36165
rect 28629 36125 28641 36159
rect 28675 36156 28687 36159
rect 28810 36156 28816 36168
rect 28675 36128 28816 36156
rect 28675 36125 28687 36128
rect 28629 36119 28687 36125
rect 28810 36116 28816 36128
rect 28868 36116 28874 36168
rect 22097 36091 22155 36097
rect 22097 36088 22109 36091
rect 20732 36060 22109 36088
rect 22097 36057 22109 36060
rect 22143 36088 22155 36091
rect 22554 36088 22560 36100
rect 22143 36060 22560 36088
rect 22143 36057 22155 36060
rect 22097 36051 22155 36057
rect 22554 36048 22560 36060
rect 22612 36048 22618 36100
rect 22922 36048 22928 36100
rect 22980 36088 22986 36100
rect 25498 36088 25504 36100
rect 22980 36060 25504 36088
rect 22980 36048 22986 36060
rect 25498 36048 25504 36060
rect 25556 36088 25562 36100
rect 27890 36088 27896 36100
rect 25556 36060 27896 36088
rect 25556 36048 25562 36060
rect 27890 36048 27896 36060
rect 27948 36048 27954 36100
rect 11606 36020 11612 36032
rect 11567 35992 11612 36020
rect 11606 35980 11612 35992
rect 11664 35980 11670 36032
rect 20809 36023 20867 36029
rect 20809 35989 20821 36023
rect 20855 36020 20867 36023
rect 21358 36020 21364 36032
rect 20855 35992 21364 36020
rect 20855 35989 20867 35992
rect 20809 35983 20867 35989
rect 21358 35980 21364 35992
rect 21416 35980 21422 36032
rect 22186 35980 22192 36032
rect 22244 36020 22250 36032
rect 22297 36023 22355 36029
rect 22297 36020 22309 36023
rect 22244 35992 22309 36020
rect 22244 35980 22250 35992
rect 22297 35989 22309 35992
rect 22343 35989 22355 36023
rect 22462 36020 22468 36032
rect 22423 35992 22468 36020
rect 22297 35983 22355 35989
rect 22462 35980 22468 35992
rect 22520 35980 22526 36032
rect 25682 35980 25688 36032
rect 25740 36029 25746 36032
rect 25740 36023 25759 36029
rect 25747 35989 25759 36023
rect 25866 36020 25872 36032
rect 25827 35992 25872 36020
rect 25740 35983 25759 35989
rect 25740 35980 25746 35983
rect 25866 35980 25872 35992
rect 25924 35980 25930 36032
rect 25958 35980 25964 36032
rect 26016 36020 26022 36032
rect 28534 36020 28540 36032
rect 26016 35992 28540 36020
rect 26016 35980 26022 35992
rect 28534 35980 28540 35992
rect 28592 35980 28598 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 12986 35776 12992 35828
rect 13044 35816 13050 35828
rect 13541 35819 13599 35825
rect 13541 35816 13553 35819
rect 13044 35788 13553 35816
rect 13044 35776 13050 35788
rect 13541 35785 13553 35788
rect 13587 35785 13599 35819
rect 13541 35779 13599 35785
rect 14274 35776 14280 35828
rect 14332 35816 14338 35828
rect 15102 35816 15108 35828
rect 14332 35788 15108 35816
rect 14332 35776 14338 35788
rect 15102 35776 15108 35788
rect 15160 35776 15166 35828
rect 15746 35776 15752 35828
rect 15804 35816 15810 35828
rect 16666 35816 16672 35828
rect 15804 35788 16672 35816
rect 15804 35776 15810 35788
rect 16666 35776 16672 35788
rect 16724 35776 16730 35828
rect 17126 35776 17132 35828
rect 17184 35816 17190 35828
rect 26053 35819 26111 35825
rect 17184 35788 26004 35816
rect 17184 35776 17190 35788
rect 10045 35751 10103 35757
rect 10045 35717 10057 35751
rect 10091 35748 10103 35751
rect 10318 35748 10324 35760
rect 10091 35720 10324 35748
rect 10091 35717 10103 35720
rect 10045 35711 10103 35717
rect 10318 35708 10324 35720
rect 10376 35708 10382 35760
rect 12434 35748 12440 35760
rect 11532 35720 12440 35748
rect 9861 35683 9919 35689
rect 9861 35649 9873 35683
rect 9907 35680 9919 35683
rect 10962 35680 10968 35692
rect 9907 35652 10968 35680
rect 9907 35649 9919 35652
rect 9861 35643 9919 35649
rect 10962 35640 10968 35652
rect 11020 35640 11026 35692
rect 11532 35689 11560 35720
rect 12434 35708 12440 35720
rect 12492 35708 12498 35760
rect 12894 35708 12900 35760
rect 12952 35748 12958 35760
rect 16936 35751 16994 35757
rect 12952 35720 16804 35748
rect 12952 35708 12958 35720
rect 11517 35683 11575 35689
rect 11517 35649 11529 35683
rect 11563 35649 11575 35683
rect 11517 35643 11575 35649
rect 11606 35640 11612 35692
rect 11664 35680 11670 35692
rect 13372 35689 13400 35720
rect 11773 35683 11831 35689
rect 11773 35680 11785 35683
rect 11664 35652 11785 35680
rect 11664 35640 11670 35652
rect 11773 35649 11785 35652
rect 11819 35649 11831 35683
rect 11773 35643 11831 35649
rect 13357 35683 13415 35689
rect 13357 35649 13369 35683
rect 13403 35649 13415 35683
rect 15470 35680 15476 35692
rect 15431 35652 15476 35680
rect 13357 35643 13415 35649
rect 15470 35640 15476 35652
rect 15528 35640 15534 35692
rect 15565 35683 15623 35689
rect 15565 35649 15577 35683
rect 15611 35649 15623 35683
rect 15746 35680 15752 35692
rect 15707 35652 15752 35680
rect 15565 35643 15623 35649
rect 12986 35572 12992 35624
rect 13044 35612 13050 35624
rect 15580 35612 15608 35643
rect 15746 35640 15752 35652
rect 15804 35640 15810 35692
rect 15838 35640 15844 35692
rect 15896 35680 15902 35692
rect 16666 35680 16672 35692
rect 15896 35652 15941 35680
rect 16627 35652 16672 35680
rect 15896 35640 15902 35652
rect 16666 35640 16672 35652
rect 16724 35640 16730 35692
rect 16776 35680 16804 35720
rect 16936 35717 16948 35751
rect 16982 35748 16994 35751
rect 21910 35748 21916 35760
rect 16982 35720 21916 35748
rect 16982 35717 16994 35720
rect 16936 35711 16994 35717
rect 21910 35708 21916 35720
rect 21968 35708 21974 35760
rect 22281 35751 22339 35757
rect 22281 35717 22293 35751
rect 22327 35748 22339 35751
rect 22738 35748 22744 35760
rect 22327 35720 22744 35748
rect 22327 35717 22339 35720
rect 22281 35711 22339 35717
rect 22738 35708 22744 35720
rect 22796 35708 22802 35760
rect 25038 35748 25044 35760
rect 23124 35720 25044 35748
rect 19061 35683 19119 35689
rect 19061 35680 19073 35683
rect 16776 35652 19073 35680
rect 19061 35649 19073 35652
rect 19107 35649 19119 35683
rect 19061 35643 19119 35649
rect 19150 35640 19156 35692
rect 19208 35680 19214 35692
rect 19889 35683 19947 35689
rect 19208 35652 19840 35680
rect 19208 35640 19214 35652
rect 19702 35612 19708 35624
rect 13044 35584 15608 35612
rect 19663 35584 19708 35612
rect 13044 35572 13050 35584
rect 19702 35572 19708 35584
rect 19760 35572 19766 35624
rect 19812 35612 19840 35652
rect 19889 35649 19901 35683
rect 19935 35680 19947 35683
rect 20070 35680 20076 35692
rect 19935 35652 20076 35680
rect 19935 35649 19947 35652
rect 19889 35643 19947 35649
rect 20070 35640 20076 35652
rect 20128 35640 20134 35692
rect 20533 35683 20591 35689
rect 20533 35680 20545 35683
rect 20180 35652 20545 35680
rect 20180 35612 20208 35652
rect 20533 35649 20545 35652
rect 20579 35649 20591 35683
rect 20533 35643 20591 35649
rect 20717 35683 20775 35689
rect 20717 35649 20729 35683
rect 20763 35680 20775 35683
rect 21450 35680 21456 35692
rect 20763 35652 21456 35680
rect 20763 35649 20775 35652
rect 20717 35643 20775 35649
rect 21450 35640 21456 35652
rect 21508 35640 21514 35692
rect 22922 35680 22928 35692
rect 21560 35652 22928 35680
rect 20622 35612 20628 35624
rect 19812 35584 20208 35612
rect 20583 35584 20628 35612
rect 20622 35572 20628 35584
rect 20680 35572 20686 35624
rect 15470 35504 15476 35556
rect 15528 35544 15534 35556
rect 15654 35544 15660 35556
rect 15528 35516 15660 35544
rect 15528 35504 15534 35516
rect 15654 35504 15660 35516
rect 15712 35504 15718 35556
rect 19245 35547 19303 35553
rect 19245 35513 19257 35547
rect 19291 35544 19303 35547
rect 21560 35544 21588 35652
rect 22922 35640 22928 35652
rect 22980 35640 22986 35692
rect 23124 35689 23152 35720
rect 25038 35708 25044 35720
rect 25096 35708 25102 35760
rect 25774 35708 25780 35760
rect 25832 35748 25838 35760
rect 25869 35751 25927 35757
rect 25869 35748 25881 35751
rect 25832 35720 25881 35748
rect 25832 35708 25838 35720
rect 25869 35717 25881 35720
rect 25915 35717 25927 35751
rect 25869 35711 25927 35717
rect 23109 35683 23167 35689
rect 23109 35649 23121 35683
rect 23155 35649 23167 35683
rect 23109 35643 23167 35649
rect 23376 35683 23434 35689
rect 23376 35649 23388 35683
rect 23422 35680 23434 35683
rect 24302 35680 24308 35692
rect 23422 35652 24308 35680
rect 23422 35649 23434 35652
rect 23376 35643 23434 35649
rect 24302 35640 24308 35652
rect 24360 35640 24366 35692
rect 25976 35680 26004 35788
rect 26053 35785 26065 35819
rect 26099 35816 26111 35819
rect 26510 35816 26516 35828
rect 26099 35788 26516 35816
rect 26099 35785 26111 35788
rect 26053 35779 26111 35785
rect 26510 35776 26516 35788
rect 26568 35776 26574 35828
rect 28103 35819 28161 35825
rect 28103 35785 28115 35819
rect 28149 35816 28161 35819
rect 28258 35816 28264 35828
rect 28149 35788 28264 35816
rect 28149 35785 28161 35788
rect 28103 35779 28161 35785
rect 28258 35776 28264 35788
rect 28316 35776 28322 35828
rect 28626 35776 28632 35828
rect 28684 35816 28690 35828
rect 28813 35819 28871 35825
rect 28813 35816 28825 35819
rect 28684 35788 28825 35816
rect 28684 35776 28690 35788
rect 28813 35785 28825 35788
rect 28859 35785 28871 35819
rect 28813 35779 28871 35785
rect 29733 35819 29791 35825
rect 29733 35785 29745 35819
rect 29779 35785 29791 35819
rect 29733 35779 29791 35785
rect 27890 35748 27896 35760
rect 27851 35720 27896 35748
rect 27890 35708 27896 35720
rect 27948 35708 27954 35760
rect 29748 35748 29776 35779
rect 30377 35751 30435 35757
rect 30377 35748 30389 35751
rect 28184 35720 29776 35748
rect 29840 35720 30389 35748
rect 28184 35680 28212 35720
rect 25976 35652 28212 35680
rect 28442 35640 28448 35692
rect 28500 35680 28506 35692
rect 28718 35680 28724 35692
rect 28500 35652 28724 35680
rect 28500 35640 28506 35652
rect 28718 35640 28724 35652
rect 28776 35640 28782 35692
rect 28810 35640 28816 35692
rect 28868 35680 28874 35692
rect 28905 35683 28963 35689
rect 28905 35680 28917 35683
rect 28868 35652 28917 35680
rect 28868 35640 28874 35652
rect 28905 35649 28917 35652
rect 28951 35649 28963 35683
rect 28905 35643 28963 35649
rect 29549 35683 29607 35689
rect 29549 35649 29561 35683
rect 29595 35680 29607 35683
rect 29730 35680 29736 35692
rect 29595 35652 29736 35680
rect 29595 35649 29607 35652
rect 29549 35643 29607 35649
rect 29730 35640 29736 35652
rect 29788 35640 29794 35692
rect 22462 35572 22468 35624
rect 22520 35572 22526 35624
rect 28092 35584 28488 35612
rect 19291 35516 21588 35544
rect 19291 35513 19303 35516
rect 19245 35507 19303 35513
rect 21634 35504 21640 35556
rect 21692 35544 21698 35556
rect 21913 35547 21971 35553
rect 21913 35544 21925 35547
rect 21692 35516 21925 35544
rect 21692 35504 21698 35516
rect 21913 35513 21925 35516
rect 21959 35513 21971 35547
rect 22480 35544 22508 35572
rect 25498 35544 25504 35556
rect 21913 35507 21971 35513
rect 22296 35516 22508 35544
rect 25459 35516 25504 35544
rect 9950 35436 9956 35488
rect 10008 35476 10014 35488
rect 10229 35479 10287 35485
rect 10229 35476 10241 35479
rect 10008 35448 10241 35476
rect 10008 35436 10014 35448
rect 10229 35445 10241 35448
rect 10275 35445 10287 35479
rect 10229 35439 10287 35445
rect 12250 35436 12256 35488
rect 12308 35476 12314 35488
rect 12897 35479 12955 35485
rect 12897 35476 12909 35479
rect 12308 35448 12909 35476
rect 12308 35436 12314 35448
rect 12897 35445 12909 35448
rect 12943 35445 12955 35479
rect 12897 35439 12955 35445
rect 13998 35436 14004 35488
rect 14056 35476 14062 35488
rect 15289 35479 15347 35485
rect 15289 35476 15301 35479
rect 14056 35448 15301 35476
rect 14056 35436 14062 35448
rect 15289 35445 15301 35448
rect 15335 35445 15347 35479
rect 15289 35439 15347 35445
rect 16942 35436 16948 35488
rect 17000 35476 17006 35488
rect 18049 35479 18107 35485
rect 18049 35476 18061 35479
rect 17000 35448 18061 35476
rect 17000 35436 17006 35448
rect 18049 35445 18061 35448
rect 18095 35445 18107 35479
rect 18049 35439 18107 35445
rect 20073 35479 20131 35485
rect 20073 35445 20085 35479
rect 20119 35476 20131 35479
rect 20990 35476 20996 35488
rect 20119 35448 20996 35476
rect 20119 35445 20131 35448
rect 20073 35439 20131 35445
rect 20990 35436 20996 35448
rect 21048 35436 21054 35488
rect 22296 35485 22324 35516
rect 25498 35504 25504 35516
rect 25556 35504 25562 35556
rect 22281 35479 22339 35485
rect 22281 35445 22293 35479
rect 22327 35445 22339 35479
rect 22462 35476 22468 35488
rect 22423 35448 22468 35476
rect 22281 35439 22339 35445
rect 22462 35436 22468 35448
rect 22520 35436 22526 35488
rect 24486 35476 24492 35488
rect 24447 35448 24492 35476
rect 24486 35436 24492 35448
rect 24544 35436 24550 35488
rect 25866 35476 25872 35488
rect 25827 35448 25872 35476
rect 25866 35436 25872 35448
rect 25924 35436 25930 35488
rect 28092 35485 28120 35584
rect 28166 35504 28172 35556
rect 28224 35504 28230 35556
rect 28077 35479 28135 35485
rect 28077 35445 28089 35479
rect 28123 35445 28135 35479
rect 28184 35476 28212 35504
rect 28261 35479 28319 35485
rect 28261 35476 28273 35479
rect 28184 35448 28273 35476
rect 28077 35439 28135 35445
rect 28261 35445 28273 35448
rect 28307 35445 28319 35479
rect 28460 35476 28488 35584
rect 28534 35504 28540 35556
rect 28592 35544 28598 35556
rect 29840 35544 29868 35720
rect 30377 35717 30389 35720
rect 30423 35717 30435 35751
rect 30377 35711 30435 35717
rect 30392 35680 30420 35711
rect 30558 35708 30564 35760
rect 30616 35757 30622 35760
rect 30616 35751 30635 35757
rect 30623 35717 30635 35751
rect 30616 35711 30635 35717
rect 30616 35708 30622 35711
rect 30834 35680 30840 35692
rect 30392 35652 30840 35680
rect 30834 35640 30840 35652
rect 30892 35640 30898 35692
rect 37550 35612 37556 35624
rect 28592 35516 29868 35544
rect 29932 35584 37556 35612
rect 28592 35504 28598 35516
rect 29932 35476 29960 35584
rect 37550 35572 37556 35584
rect 37608 35572 37614 35624
rect 32122 35544 32128 35556
rect 30576 35516 32128 35544
rect 30576 35485 30604 35516
rect 32122 35504 32128 35516
rect 32180 35504 32186 35556
rect 28460 35448 29960 35476
rect 30561 35479 30619 35485
rect 28261 35439 28319 35445
rect 30561 35445 30573 35479
rect 30607 35445 30619 35479
rect 30742 35476 30748 35488
rect 30703 35448 30748 35476
rect 30561 35439 30619 35445
rect 30742 35436 30748 35448
rect 30800 35436 30806 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 9858 35272 9864 35284
rect 9819 35244 9864 35272
rect 9858 35232 9864 35244
rect 9916 35232 9922 35284
rect 11790 35272 11796 35284
rect 11751 35244 11796 35272
rect 11790 35232 11796 35244
rect 11848 35232 11854 35284
rect 14090 35272 14096 35284
rect 11992 35244 14096 35272
rect 9858 35096 9864 35148
rect 9916 35136 9922 35148
rect 11333 35139 11391 35145
rect 11333 35136 11345 35139
rect 9916 35108 10272 35136
rect 9916 35096 9922 35108
rect 10244 35077 10272 35108
rect 10336 35108 11345 35136
rect 10336 35077 10364 35108
rect 11333 35105 11345 35108
rect 11379 35105 11391 35139
rect 11333 35099 11391 35105
rect 10137 35071 10195 35077
rect 10137 35037 10149 35071
rect 10183 35037 10195 35071
rect 10137 35031 10195 35037
rect 10229 35071 10287 35077
rect 10229 35037 10241 35071
rect 10275 35037 10287 35071
rect 10229 35031 10287 35037
rect 10321 35071 10379 35077
rect 10321 35037 10333 35071
rect 10367 35037 10379 35071
rect 10502 35068 10508 35080
rect 10463 35040 10508 35068
rect 10321 35031 10379 35037
rect 10152 34932 10180 35031
rect 10502 35028 10508 35040
rect 10560 35028 10566 35080
rect 10962 35068 10968 35080
rect 10923 35040 10968 35068
rect 10962 35028 10968 35040
rect 11020 35028 11026 35080
rect 11146 35068 11152 35080
rect 11107 35040 11152 35068
rect 11146 35028 11152 35040
rect 11204 35028 11210 35080
rect 11992 35077 12020 35244
rect 14090 35232 14096 35244
rect 14148 35272 14154 35284
rect 14148 35244 15516 35272
rect 14148 35232 14154 35244
rect 12710 35204 12716 35216
rect 12671 35176 12716 35204
rect 12710 35164 12716 35176
rect 12768 35164 12774 35216
rect 14458 35164 14464 35216
rect 14516 35204 14522 35216
rect 15488 35204 15516 35244
rect 15746 35232 15752 35284
rect 15804 35272 15810 35284
rect 16761 35275 16819 35281
rect 16761 35272 16773 35275
rect 15804 35244 16773 35272
rect 15804 35232 15810 35244
rect 16761 35241 16773 35244
rect 16807 35241 16819 35275
rect 17954 35272 17960 35284
rect 17915 35244 17960 35272
rect 16761 35235 16819 35241
rect 17954 35232 17960 35244
rect 18012 35232 18018 35284
rect 19242 35272 19248 35284
rect 19203 35244 19248 35272
rect 19242 35232 19248 35244
rect 19300 35232 19306 35284
rect 21726 35232 21732 35284
rect 21784 35272 21790 35284
rect 21821 35275 21879 35281
rect 21821 35272 21833 35275
rect 21784 35244 21833 35272
rect 21784 35232 21790 35244
rect 21821 35241 21833 35244
rect 21867 35241 21879 35275
rect 21821 35235 21879 35241
rect 21910 35232 21916 35284
rect 21968 35272 21974 35284
rect 22281 35275 22339 35281
rect 22281 35272 22293 35275
rect 21968 35244 22293 35272
rect 21968 35232 21974 35244
rect 22281 35241 22293 35244
rect 22327 35241 22339 35275
rect 22281 35235 22339 35241
rect 23661 35275 23719 35281
rect 23661 35241 23673 35275
rect 23707 35241 23719 35275
rect 28166 35272 28172 35284
rect 28127 35244 28172 35272
rect 23661 35235 23719 35241
rect 14516 35176 15424 35204
rect 15488 35176 15783 35204
rect 14516 35164 14522 35176
rect 15289 35139 15347 35145
rect 15289 35136 15301 35139
rect 14108 35108 15301 35136
rect 11793 35071 11851 35077
rect 11793 35037 11805 35071
rect 11839 35037 11851 35071
rect 11793 35031 11851 35037
rect 11977 35071 12035 35077
rect 11977 35037 11989 35071
rect 12023 35037 12035 35071
rect 11977 35031 12035 35037
rect 12529 35071 12587 35077
rect 12529 35037 12541 35071
rect 12575 35068 12587 35071
rect 12894 35068 12900 35080
rect 12575 35040 12900 35068
rect 12575 35037 12587 35040
rect 12529 35031 12587 35037
rect 11808 35000 11836 35031
rect 12894 35028 12900 35040
rect 12952 35068 12958 35080
rect 13170 35068 13176 35080
rect 12952 35040 13176 35068
rect 12952 35028 12958 35040
rect 13170 35028 13176 35040
rect 13228 35028 13234 35080
rect 14108 35077 14136 35108
rect 15289 35105 15301 35108
rect 15335 35105 15347 35139
rect 15396 35136 15424 35176
rect 15396 35108 15700 35136
rect 15289 35099 15347 35105
rect 14093 35071 14151 35077
rect 14093 35037 14105 35071
rect 14139 35037 14151 35071
rect 14093 35031 14151 35037
rect 14182 35028 14188 35080
rect 14240 35068 14246 35080
rect 14642 35077 14648 35080
rect 14599 35071 14648 35077
rect 14240 35040 14285 35068
rect 14240 35028 14246 35040
rect 14599 35037 14611 35071
rect 14645 35037 14648 35071
rect 14599 35031 14648 35037
rect 14642 35028 14648 35031
rect 14700 35028 14706 35080
rect 15378 35028 15384 35080
rect 15436 35068 15442 35080
rect 15672 35077 15700 35108
rect 15473 35071 15531 35077
rect 15473 35068 15485 35071
rect 15436 35040 15485 35068
rect 15436 35028 15442 35040
rect 15473 35037 15485 35040
rect 15519 35037 15531 35071
rect 15473 35031 15531 35037
rect 15657 35071 15715 35077
rect 15657 35037 15669 35071
rect 15703 35037 15715 35071
rect 15755 35068 15783 35176
rect 16482 35164 16488 35216
rect 16540 35204 16546 35216
rect 21634 35204 21640 35216
rect 16540 35176 19380 35204
rect 21595 35176 21640 35204
rect 16540 35164 16546 35176
rect 15933 35139 15991 35145
rect 15933 35105 15945 35139
rect 15979 35136 15991 35139
rect 16206 35136 16212 35148
rect 15979 35108 16212 35136
rect 15979 35105 15991 35108
rect 15933 35099 15991 35105
rect 16206 35096 16212 35108
rect 16264 35136 16270 35148
rect 19150 35136 19156 35148
rect 16264 35108 19156 35136
rect 16264 35096 16270 35108
rect 19150 35096 19156 35108
rect 19208 35096 19214 35148
rect 16393 35071 16451 35077
rect 16393 35068 16405 35071
rect 15755 35040 16405 35068
rect 15657 35031 15715 35037
rect 16393 35037 16405 35040
rect 16439 35037 16451 35071
rect 16393 35031 16451 35037
rect 16577 35071 16635 35077
rect 16577 35037 16589 35071
rect 16623 35068 16635 35071
rect 17678 35068 17684 35080
rect 16623 35040 17684 35068
rect 16623 35037 16635 35040
rect 16577 35031 16635 35037
rect 17678 35028 17684 35040
rect 17736 35028 17742 35080
rect 17957 35071 18015 35077
rect 17957 35037 17969 35071
rect 18003 35037 18015 35071
rect 17957 35031 18015 35037
rect 18141 35071 18199 35077
rect 18141 35037 18153 35071
rect 18187 35068 18199 35071
rect 18414 35068 18420 35080
rect 18187 35040 18420 35068
rect 18187 35037 18199 35040
rect 18141 35031 18199 35037
rect 12434 35000 12440 35012
rect 11808 34972 12440 35000
rect 12434 34960 12440 34972
rect 12492 34960 12498 35012
rect 12986 35000 12992 35012
rect 12544 34972 12992 35000
rect 12544 34932 12572 34972
rect 12986 34960 12992 34972
rect 13044 34960 13050 35012
rect 14366 35000 14372 35012
rect 14327 34972 14372 35000
rect 14366 34960 14372 34972
rect 14424 34960 14430 35012
rect 14461 35003 14519 35009
rect 14461 34969 14473 35003
rect 14507 35000 14519 35003
rect 14918 35000 14924 35012
rect 14507 34972 14924 35000
rect 14507 34969 14519 34972
rect 14461 34963 14519 34969
rect 14918 34960 14924 34972
rect 14976 34960 14982 35012
rect 15565 35003 15623 35009
rect 15565 34969 15577 35003
rect 15611 35000 15623 35003
rect 15795 35003 15853 35009
rect 15611 34972 15700 35000
rect 15611 34969 15623 34972
rect 15565 34963 15623 34969
rect 15672 34944 15700 34972
rect 15795 34969 15807 35003
rect 15841 35000 15853 35003
rect 17972 35000 18000 35031
rect 18414 35028 18420 35040
rect 18472 35028 18478 35080
rect 19245 35071 19303 35077
rect 19245 35068 19257 35071
rect 19168 35040 19257 35068
rect 19168 35012 19196 35040
rect 19245 35037 19257 35040
rect 19291 35037 19303 35071
rect 19245 35031 19303 35037
rect 18874 35000 18880 35012
rect 15841 34972 18880 35000
rect 15841 34969 15853 34972
rect 15795 34963 15853 34969
rect 18874 34960 18880 34972
rect 18932 34960 18938 35012
rect 19150 34960 19156 35012
rect 19208 34960 19214 35012
rect 10152 34904 12572 34932
rect 14550 34892 14556 34944
rect 14608 34932 14614 34944
rect 14737 34935 14795 34941
rect 14737 34932 14749 34935
rect 14608 34904 14749 34932
rect 14608 34892 14614 34904
rect 14737 34901 14749 34904
rect 14783 34901 14795 34935
rect 14737 34895 14795 34901
rect 15654 34892 15660 34944
rect 15712 34892 15718 34944
rect 19352 34932 19380 35176
rect 21634 35164 21640 35176
rect 21692 35164 21698 35216
rect 19702 35096 19708 35148
rect 19760 35136 19766 35148
rect 22186 35136 22192 35148
rect 19760 35108 20668 35136
rect 19760 35096 19766 35108
rect 20640 35080 20668 35108
rect 21376 35108 22192 35136
rect 19429 35071 19487 35077
rect 19429 35037 19441 35071
rect 19475 35068 19487 35071
rect 20346 35068 20352 35080
rect 19475 35040 20352 35068
rect 19475 35037 19487 35040
rect 19429 35031 19487 35037
rect 20346 35028 20352 35040
rect 20404 35028 20410 35080
rect 20622 35028 20628 35080
rect 20680 35068 20686 35080
rect 20717 35071 20775 35077
rect 20717 35068 20729 35071
rect 20680 35040 20729 35068
rect 20680 35028 20686 35040
rect 20717 35037 20729 35040
rect 20763 35037 20775 35071
rect 20717 35031 20775 35037
rect 20901 35071 20959 35077
rect 20901 35037 20913 35071
rect 20947 35068 20959 35071
rect 20990 35068 20996 35080
rect 20947 35040 20996 35068
rect 20947 35037 20959 35040
rect 20901 35031 20959 35037
rect 20990 35028 20996 35040
rect 21048 35028 21054 35080
rect 21376 35009 21404 35108
rect 22186 35096 22192 35108
rect 22244 35096 22250 35148
rect 23676 35136 23704 35235
rect 28166 35232 28172 35244
rect 28224 35232 28230 35284
rect 30374 35272 30380 35284
rect 30335 35244 30380 35272
rect 30374 35232 30380 35244
rect 30432 35232 30438 35284
rect 31018 35272 31024 35284
rect 30979 35244 31024 35272
rect 31018 35232 31024 35244
rect 31076 35232 31082 35284
rect 25409 35207 25467 35213
rect 25409 35173 25421 35207
rect 25455 35204 25467 35207
rect 25498 35204 25504 35216
rect 25455 35176 25504 35204
rect 25455 35173 25467 35176
rect 25409 35167 25467 35173
rect 25498 35164 25504 35176
rect 25556 35204 25562 35216
rect 25961 35207 26019 35213
rect 25961 35204 25973 35207
rect 25556 35176 25973 35204
rect 25556 35164 25562 35176
rect 25961 35173 25973 35176
rect 26007 35173 26019 35207
rect 30190 35204 30196 35216
rect 30151 35176 30196 35204
rect 25961 35167 26019 35173
rect 30190 35164 30196 35176
rect 30248 35164 30254 35216
rect 30466 35164 30472 35216
rect 30524 35204 30530 35216
rect 31205 35207 31263 35213
rect 31205 35204 31217 35207
rect 30524 35176 31217 35204
rect 30524 35164 30530 35176
rect 31205 35173 31217 35176
rect 31251 35173 31263 35207
rect 31205 35167 31263 35173
rect 32398 35136 32404 35148
rect 23676 35108 32404 35136
rect 32398 35096 32404 35108
rect 32456 35096 32462 35148
rect 22462 35068 22468 35080
rect 22423 35040 22468 35068
rect 22462 35028 22468 35040
rect 22520 35028 22526 35080
rect 25958 35068 25964 35080
rect 25919 35040 25964 35068
rect 25958 35028 25964 35040
rect 26016 35028 26022 35080
rect 26145 35071 26203 35077
rect 26145 35037 26157 35071
rect 26191 35068 26203 35071
rect 26326 35068 26332 35080
rect 26191 35040 26332 35068
rect 26191 35037 26203 35040
rect 26145 35031 26203 35037
rect 26326 35028 26332 35040
rect 26384 35028 26390 35080
rect 27798 35068 27804 35080
rect 27759 35040 27804 35068
rect 27798 35028 27804 35040
rect 27856 35028 27862 35080
rect 28534 35028 28540 35080
rect 28592 35068 28598 35080
rect 28813 35071 28871 35077
rect 28813 35068 28825 35071
rect 28592 35040 28825 35068
rect 28592 35028 28598 35040
rect 28813 35037 28825 35040
rect 28859 35037 28871 35071
rect 28813 35031 28871 35037
rect 28997 35071 29055 35077
rect 28997 35037 29009 35071
rect 29043 35068 29055 35071
rect 29086 35068 29092 35080
rect 29043 35040 29092 35068
rect 29043 35037 29055 35040
rect 28997 35031 29055 35037
rect 29086 35028 29092 35040
rect 29144 35028 29150 35080
rect 29917 35071 29975 35077
rect 29917 35037 29929 35071
rect 29963 35068 29975 35071
rect 30558 35068 30564 35080
rect 29963 35040 30564 35068
rect 29963 35037 29975 35040
rect 29917 35031 29975 35037
rect 30558 35028 30564 35040
rect 30616 35068 30622 35080
rect 31110 35068 31116 35080
rect 30616 35040 31116 35068
rect 30616 35028 30622 35040
rect 31110 35028 31116 35040
rect 31168 35028 31174 35080
rect 20809 35003 20867 35009
rect 20809 34969 20821 35003
rect 20855 35000 20867 35003
rect 21361 35003 21419 35009
rect 21361 35000 21373 35003
rect 20855 34972 21373 35000
rect 20855 34969 20867 34972
rect 20809 34963 20867 34969
rect 21361 34969 21373 34972
rect 21407 34969 21419 35003
rect 21361 34963 21419 34969
rect 22554 34960 22560 35012
rect 22612 35000 22618 35012
rect 23477 35003 23535 35009
rect 23477 35000 23489 35003
rect 22612 34972 23489 35000
rect 22612 34960 22618 34972
rect 23477 34969 23489 34972
rect 23523 34969 23535 35003
rect 23477 34963 23535 34969
rect 23693 35003 23751 35009
rect 23693 34969 23705 35003
rect 23739 35000 23751 35003
rect 23934 35000 23940 35012
rect 23739 34972 23940 35000
rect 23739 34969 23751 34972
rect 23693 34963 23751 34969
rect 23934 34960 23940 34972
rect 23992 34960 23998 35012
rect 25041 35003 25099 35009
rect 25041 34969 25053 35003
rect 25087 35000 25099 35003
rect 25682 35000 25688 35012
rect 25087 34972 25688 35000
rect 25087 34969 25099 34972
rect 25041 34963 25099 34969
rect 25682 34960 25688 34972
rect 25740 34960 25746 35012
rect 28169 35003 28227 35009
rect 28169 34969 28181 35003
rect 28215 35000 28227 35003
rect 28905 35003 28963 35009
rect 28905 35000 28917 35003
rect 28215 34972 28917 35000
rect 28215 34969 28227 34972
rect 28169 34963 28227 34969
rect 28905 34969 28917 34972
rect 28951 34969 28963 35003
rect 30834 35000 30840 35012
rect 30795 34972 30840 35000
rect 28905 34963 28963 34969
rect 30834 34960 30840 34972
rect 30892 34960 30898 35012
rect 23566 34932 23572 34944
rect 19352 34904 23572 34932
rect 23566 34892 23572 34904
rect 23624 34892 23630 34944
rect 23842 34932 23848 34944
rect 23803 34904 23848 34932
rect 23842 34892 23848 34904
rect 23900 34892 23906 34944
rect 25314 34892 25320 34944
rect 25372 34932 25378 34944
rect 25501 34935 25559 34941
rect 25501 34932 25513 34935
rect 25372 34904 25513 34932
rect 25372 34892 25378 34904
rect 25501 34901 25513 34904
rect 25547 34901 25559 34935
rect 25501 34895 25559 34901
rect 28074 34892 28080 34944
rect 28132 34932 28138 34944
rect 28353 34935 28411 34941
rect 28353 34932 28365 34935
rect 28132 34904 28365 34932
rect 28132 34892 28138 34904
rect 28353 34901 28365 34904
rect 28399 34901 28411 34935
rect 28353 34895 28411 34901
rect 30374 34892 30380 34944
rect 30432 34932 30438 34944
rect 31047 34935 31105 34941
rect 31047 34932 31059 34935
rect 30432 34904 31059 34932
rect 30432 34892 30438 34904
rect 31047 34901 31059 34904
rect 31093 34932 31105 34935
rect 31570 34932 31576 34944
rect 31093 34904 31576 34932
rect 31093 34901 31105 34904
rect 31047 34895 31105 34901
rect 31570 34892 31576 34904
rect 31628 34892 31634 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 8665 34731 8723 34737
rect 8665 34697 8677 34731
rect 8711 34728 8723 34731
rect 9582 34728 9588 34740
rect 8711 34700 9588 34728
rect 8711 34697 8723 34700
rect 8665 34691 8723 34697
rect 9582 34688 9588 34700
rect 9640 34688 9646 34740
rect 12618 34688 12624 34740
rect 12676 34688 12682 34740
rect 12713 34731 12771 34737
rect 12713 34697 12725 34731
rect 12759 34728 12771 34731
rect 13722 34728 13728 34740
rect 12759 34700 13728 34728
rect 12759 34697 12771 34700
rect 12713 34691 12771 34697
rect 13722 34688 13728 34700
rect 13780 34688 13786 34740
rect 13906 34688 13912 34740
rect 13964 34728 13970 34740
rect 14277 34731 14335 34737
rect 14277 34728 14289 34731
rect 13964 34700 14289 34728
rect 13964 34688 13970 34700
rect 14277 34697 14289 34700
rect 14323 34697 14335 34731
rect 17770 34728 17776 34740
rect 14277 34691 14335 34697
rect 16689 34700 17776 34728
rect 10410 34660 10416 34672
rect 9140 34632 10416 34660
rect 8938 34592 8944 34604
rect 8899 34564 8944 34592
rect 8938 34552 8944 34564
rect 8996 34552 9002 34604
rect 9140 34601 9168 34632
rect 10410 34620 10416 34632
rect 10468 34620 10474 34672
rect 12437 34663 12495 34669
rect 12437 34629 12449 34663
rect 12483 34660 12495 34663
rect 12636 34660 12664 34688
rect 12894 34660 12900 34672
rect 12483 34632 12900 34660
rect 12483 34629 12495 34632
rect 12437 34623 12495 34629
rect 12894 34620 12900 34632
rect 12952 34620 12958 34672
rect 16482 34660 16488 34672
rect 13832 34632 16488 34660
rect 9033 34595 9091 34601
rect 9033 34561 9045 34595
rect 9079 34561 9091 34595
rect 9033 34555 9091 34561
rect 9125 34595 9183 34601
rect 9125 34561 9137 34595
rect 9171 34561 9183 34595
rect 9125 34555 9183 34561
rect 9309 34595 9367 34601
rect 9309 34561 9321 34595
rect 9355 34592 9367 34595
rect 12066 34592 12072 34604
rect 9355 34564 10088 34592
rect 12027 34564 12072 34592
rect 9355 34561 9367 34564
rect 9309 34555 9367 34561
rect 9048 34524 9076 34555
rect 9766 34524 9772 34536
rect 9048 34496 9628 34524
rect 9727 34496 9772 34524
rect 9600 34456 9628 34496
rect 9766 34484 9772 34496
rect 9824 34484 9830 34536
rect 10060 34533 10088 34564
rect 12066 34552 12072 34564
rect 12124 34552 12130 34604
rect 12250 34601 12256 34604
rect 12217 34595 12256 34601
rect 12217 34561 12229 34595
rect 12217 34555 12256 34561
rect 12250 34552 12256 34555
rect 12308 34552 12314 34604
rect 12618 34601 12624 34604
rect 12345 34595 12403 34601
rect 12345 34561 12357 34595
rect 12391 34561 12403 34595
rect 12345 34555 12403 34561
rect 12575 34595 12624 34601
rect 12575 34561 12587 34595
rect 12621 34561 12624 34595
rect 12575 34555 12624 34561
rect 10045 34527 10103 34533
rect 10045 34493 10057 34527
rect 10091 34524 10103 34527
rect 10226 34524 10232 34536
rect 10091 34496 10232 34524
rect 10091 34493 10103 34496
rect 10045 34487 10103 34493
rect 10226 34484 10232 34496
rect 10284 34524 10290 34536
rect 10502 34524 10508 34536
rect 10284 34496 10508 34524
rect 10284 34484 10290 34496
rect 10502 34484 10508 34496
rect 10560 34484 10566 34536
rect 12360 34524 12388 34555
rect 12618 34552 12624 34555
rect 12676 34552 12682 34604
rect 13630 34592 13636 34604
rect 13591 34564 13636 34592
rect 13630 34552 13636 34564
rect 13688 34552 13694 34604
rect 13832 34601 13860 34632
rect 16482 34620 16488 34632
rect 16540 34620 16546 34672
rect 13781 34595 13860 34601
rect 13781 34561 13793 34595
rect 13827 34564 13860 34595
rect 13909 34595 13967 34601
rect 13827 34561 13839 34564
rect 13781 34555 13839 34561
rect 13909 34561 13921 34595
rect 13955 34561 13967 34595
rect 13909 34555 13967 34561
rect 14001 34595 14059 34601
rect 14001 34561 14013 34595
rect 14047 34561 14059 34595
rect 14001 34555 14059 34561
rect 14139 34595 14197 34601
rect 14139 34561 14151 34595
rect 14185 34592 14197 34595
rect 14642 34592 14648 34604
rect 14185 34564 14648 34592
rect 14185 34561 14197 34564
rect 14139 34555 14197 34561
rect 13924 34524 13952 34555
rect 12360 34496 13952 34524
rect 14016 34524 14044 34555
rect 14642 34552 14648 34564
rect 14700 34592 14706 34604
rect 15102 34592 15108 34604
rect 14700 34564 15108 34592
rect 14700 34552 14706 34564
rect 15102 34552 15108 34564
rect 15160 34592 15166 34604
rect 15473 34595 15531 34601
rect 15473 34592 15485 34595
rect 15160 34564 15485 34592
rect 15160 34552 15166 34564
rect 15473 34561 15485 34564
rect 15519 34561 15531 34595
rect 15473 34555 15531 34561
rect 14274 34524 14280 34536
rect 14016 34496 14280 34524
rect 9858 34456 9864 34468
rect 9600 34428 9864 34456
rect 9858 34416 9864 34428
rect 9916 34416 9922 34468
rect 13924 34456 13952 34496
rect 14274 34484 14280 34496
rect 14332 34484 14338 34536
rect 15197 34527 15255 34533
rect 15197 34493 15209 34527
rect 15243 34524 15255 34527
rect 16689 34524 16717 34700
rect 17770 34688 17776 34700
rect 17828 34688 17834 34740
rect 19334 34728 19340 34740
rect 19076 34700 19340 34728
rect 17037 34663 17095 34669
rect 17037 34629 17049 34663
rect 17083 34660 17095 34663
rect 17862 34660 17868 34672
rect 17083 34632 17868 34660
rect 17083 34629 17095 34632
rect 17037 34623 17095 34629
rect 17862 34620 17868 34632
rect 17920 34620 17926 34672
rect 17954 34620 17960 34672
rect 18012 34660 18018 34672
rect 18966 34660 18972 34672
rect 18012 34632 18972 34660
rect 18012 34620 18018 34632
rect 18966 34620 18972 34632
rect 19024 34620 19030 34672
rect 19076 34669 19104 34700
rect 19334 34688 19340 34700
rect 19392 34688 19398 34740
rect 20898 34728 20904 34740
rect 20272 34700 20904 34728
rect 19061 34663 19119 34669
rect 19061 34629 19073 34663
rect 19107 34629 19119 34663
rect 19061 34623 19119 34629
rect 19150 34620 19156 34672
rect 19208 34669 19214 34672
rect 19208 34663 19237 34669
rect 19225 34629 19237 34663
rect 19208 34623 19237 34629
rect 19208 34620 19214 34623
rect 19702 34620 19708 34672
rect 19760 34660 19766 34672
rect 20165 34663 20223 34669
rect 20165 34660 20177 34663
rect 19760 34632 20177 34660
rect 19760 34620 19766 34632
rect 20165 34629 20177 34632
rect 20211 34629 20223 34663
rect 20165 34623 20223 34629
rect 16850 34592 16856 34604
rect 16811 34564 16856 34592
rect 16850 34552 16856 34564
rect 16908 34552 16914 34604
rect 16945 34595 17003 34601
rect 16945 34561 16957 34595
rect 16991 34561 17003 34595
rect 16945 34555 17003 34561
rect 15243 34496 16717 34524
rect 15243 34493 15255 34496
rect 15197 34487 15255 34493
rect 14366 34456 14372 34468
rect 13924 34428 14372 34456
rect 14366 34416 14372 34428
rect 14424 34416 14430 34468
rect 16960 34456 16988 34555
rect 17126 34552 17132 34604
rect 17184 34601 17190 34604
rect 17184 34595 17213 34601
rect 17201 34561 17213 34595
rect 17184 34555 17213 34561
rect 17313 34595 17371 34601
rect 17313 34561 17325 34595
rect 17359 34592 17371 34595
rect 18322 34592 18328 34604
rect 17359 34564 18328 34592
rect 17359 34561 17371 34564
rect 17313 34555 17371 34561
rect 17184 34552 17190 34555
rect 18322 34552 18328 34564
rect 18380 34552 18386 34604
rect 20272 34601 20300 34700
rect 20898 34688 20904 34700
rect 20956 34688 20962 34740
rect 21177 34731 21235 34737
rect 21177 34697 21189 34731
rect 21223 34728 21235 34731
rect 21634 34728 21640 34740
rect 21223 34700 21640 34728
rect 21223 34697 21235 34700
rect 21177 34691 21235 34697
rect 21634 34688 21640 34700
rect 21692 34688 21698 34740
rect 22094 34688 22100 34740
rect 22152 34728 22158 34740
rect 22189 34731 22247 34737
rect 22189 34728 22201 34731
rect 22152 34700 22201 34728
rect 22152 34688 22158 34700
rect 22189 34697 22201 34700
rect 22235 34697 22247 34731
rect 22738 34728 22744 34740
rect 22699 34700 22744 34728
rect 22189 34691 22247 34697
rect 22738 34688 22744 34700
rect 22796 34688 22802 34740
rect 23845 34731 23903 34737
rect 23845 34697 23857 34731
rect 23891 34728 23903 34731
rect 24210 34728 24216 34740
rect 23891 34700 24216 34728
rect 23891 34697 23903 34700
rect 23845 34691 23903 34697
rect 24210 34688 24216 34700
rect 24268 34688 24274 34740
rect 25774 34728 25780 34740
rect 25735 34700 25780 34728
rect 25774 34688 25780 34700
rect 25832 34688 25838 34740
rect 27982 34728 27988 34740
rect 27943 34700 27988 34728
rect 27982 34688 27988 34700
rect 28040 34688 28046 34740
rect 29730 34728 29736 34740
rect 29691 34700 29736 34728
rect 29730 34688 29736 34700
rect 29788 34688 29794 34740
rect 31573 34731 31631 34737
rect 31573 34697 31585 34731
rect 31619 34697 31631 34731
rect 31573 34691 31631 34697
rect 20346 34620 20352 34672
rect 20404 34669 20410 34672
rect 20404 34663 20453 34669
rect 20404 34629 20407 34663
rect 20441 34660 20453 34663
rect 21450 34660 21456 34672
rect 20441 34632 21456 34660
rect 20441 34629 20453 34632
rect 20404 34623 20453 34629
rect 20404 34620 20410 34623
rect 21450 34620 21456 34632
rect 21508 34620 21514 34672
rect 21818 34620 21824 34672
rect 21876 34660 21882 34672
rect 21876 34632 22692 34660
rect 21876 34620 21882 34632
rect 18877 34595 18935 34601
rect 18877 34592 18889 34595
rect 18432 34564 18889 34592
rect 17954 34456 17960 34468
rect 16960 34428 17960 34456
rect 17954 34416 17960 34428
rect 18012 34416 18018 34468
rect 16666 34388 16672 34400
rect 16627 34360 16672 34388
rect 16666 34348 16672 34360
rect 16724 34348 16730 34400
rect 16850 34348 16856 34400
rect 16908 34388 16914 34400
rect 18432 34388 18460 34564
rect 18877 34561 18889 34564
rect 18923 34561 18935 34595
rect 20073 34595 20131 34601
rect 20073 34592 20085 34595
rect 18877 34555 18935 34561
rect 19260 34564 20085 34592
rect 18892 34524 18920 34555
rect 19260 34524 19288 34564
rect 20073 34561 20085 34564
rect 20119 34561 20131 34595
rect 20073 34555 20131 34561
rect 20257 34595 20315 34601
rect 20257 34561 20269 34595
rect 20303 34561 20315 34595
rect 20257 34555 20315 34561
rect 21085 34595 21143 34601
rect 21085 34561 21097 34595
rect 21131 34561 21143 34595
rect 21085 34555 21143 34561
rect 21269 34595 21327 34601
rect 21269 34561 21281 34595
rect 21315 34592 21327 34595
rect 22005 34595 22063 34601
rect 21315 34564 21956 34592
rect 21315 34561 21327 34564
rect 21269 34555 21327 34561
rect 18892 34496 19288 34524
rect 19334 34484 19340 34536
rect 19392 34524 19398 34536
rect 20346 34524 20352 34536
rect 19392 34496 20352 34524
rect 19392 34484 19398 34496
rect 20346 34484 20352 34496
rect 20404 34484 20410 34536
rect 20533 34527 20591 34533
rect 20533 34493 20545 34527
rect 20579 34493 20591 34527
rect 21100 34524 21128 34555
rect 21818 34524 21824 34536
rect 21100 34496 21824 34524
rect 20533 34487 20591 34493
rect 18966 34416 18972 34468
rect 19024 34456 19030 34468
rect 19702 34456 19708 34468
rect 19024 34428 19708 34456
rect 19024 34416 19030 34428
rect 19702 34416 19708 34428
rect 19760 34416 19766 34468
rect 20548 34456 20576 34487
rect 21818 34484 21824 34496
rect 21876 34484 21882 34536
rect 21928 34524 21956 34564
rect 22005 34561 22017 34595
rect 22051 34592 22063 34595
rect 22094 34592 22100 34604
rect 22051 34564 22100 34592
rect 22051 34561 22063 34564
rect 22005 34555 22063 34561
rect 22094 34552 22100 34564
rect 22152 34552 22158 34604
rect 22664 34601 22692 34632
rect 23566 34620 23572 34672
rect 23624 34660 23630 34672
rect 31588 34660 31616 34691
rect 23624 34632 31616 34660
rect 23624 34620 23630 34632
rect 22649 34595 22707 34601
rect 22649 34561 22661 34595
rect 22695 34561 22707 34595
rect 22808 34595 22866 34601
rect 22808 34592 22820 34595
rect 22649 34555 22707 34561
rect 22747 34564 22820 34592
rect 22747 34524 22775 34564
rect 22808 34561 22820 34564
rect 22854 34561 22866 34595
rect 22808 34555 22866 34561
rect 25685 34595 25743 34601
rect 25685 34561 25697 34595
rect 25731 34561 25743 34595
rect 25685 34555 25743 34561
rect 25869 34595 25927 34601
rect 25869 34561 25881 34595
rect 25915 34592 25927 34595
rect 26326 34592 26332 34604
rect 25915 34564 26332 34592
rect 25915 34561 25927 34564
rect 25869 34555 25927 34561
rect 21928 34496 22775 34524
rect 20898 34456 20904 34468
rect 20548 34428 20904 34456
rect 20898 34416 20904 34428
rect 20956 34456 20962 34468
rect 22094 34456 22100 34468
rect 20956 34428 22100 34456
rect 20956 34416 20962 34428
rect 22094 34416 22100 34428
rect 22152 34416 22158 34468
rect 22747 34456 22775 34496
rect 23385 34527 23443 34533
rect 23385 34493 23397 34527
rect 23431 34524 23443 34527
rect 23934 34524 23940 34536
rect 23431 34496 23940 34524
rect 23431 34493 23443 34496
rect 23385 34487 23443 34493
rect 23934 34484 23940 34496
rect 23992 34484 23998 34536
rect 25700 34524 25728 34555
rect 26326 34552 26332 34564
rect 26384 34552 26390 34604
rect 28445 34595 28503 34601
rect 28445 34561 28457 34595
rect 28491 34592 28503 34595
rect 28534 34592 28540 34604
rect 28491 34564 28540 34592
rect 28491 34561 28503 34564
rect 28445 34555 28503 34561
rect 28534 34552 28540 34564
rect 28592 34552 28598 34604
rect 28629 34595 28687 34601
rect 28629 34561 28641 34595
rect 28675 34561 28687 34595
rect 28629 34555 28687 34561
rect 25958 34524 25964 34536
rect 25700 34496 25964 34524
rect 25958 34484 25964 34496
rect 26016 34524 26022 34536
rect 26142 34524 26148 34536
rect 26016 34496 26148 34524
rect 26016 34484 26022 34496
rect 26142 34484 26148 34496
rect 26200 34484 26206 34536
rect 27525 34527 27583 34533
rect 27525 34493 27537 34527
rect 27571 34524 27583 34527
rect 28258 34524 28264 34536
rect 27571 34496 28264 34524
rect 27571 34493 27583 34496
rect 27525 34487 27583 34493
rect 28258 34484 28264 34496
rect 28316 34484 28322 34536
rect 28644 34524 28672 34555
rect 28902 34552 28908 34604
rect 28960 34592 28966 34604
rect 30193 34595 30251 34601
rect 30193 34592 30205 34595
rect 28960 34564 30205 34592
rect 28960 34552 28966 34564
rect 30193 34561 30205 34564
rect 30239 34561 30251 34595
rect 30193 34555 30251 34561
rect 30282 34552 30288 34604
rect 30340 34552 30346 34604
rect 30460 34595 30518 34601
rect 30460 34561 30472 34595
rect 30506 34592 30518 34595
rect 31202 34592 31208 34604
rect 30506 34564 31208 34592
rect 30506 34561 30518 34564
rect 30460 34555 30518 34561
rect 31202 34552 31208 34564
rect 31260 34552 31266 34604
rect 29086 34524 29092 34536
rect 28644 34496 29092 34524
rect 29086 34484 29092 34496
rect 29144 34484 29150 34536
rect 29273 34527 29331 34533
rect 29273 34493 29285 34527
rect 29319 34524 29331 34527
rect 30300 34524 30328 34552
rect 29319 34496 30328 34524
rect 29319 34493 29331 34496
rect 29273 34487 29331 34493
rect 22830 34456 22836 34468
rect 22747 34428 22836 34456
rect 22830 34416 22836 34428
rect 22888 34416 22894 34468
rect 23290 34416 23296 34468
rect 23348 34456 23354 34468
rect 23661 34459 23719 34465
rect 23661 34456 23673 34459
rect 23348 34428 23673 34456
rect 23348 34416 23354 34428
rect 23661 34425 23673 34428
rect 23707 34425 23719 34459
rect 27798 34456 27804 34468
rect 27759 34428 27804 34456
rect 23661 34419 23719 34425
rect 27798 34416 27804 34428
rect 27856 34456 27862 34468
rect 28445 34459 28503 34465
rect 28445 34456 28457 34459
rect 27856 34428 28457 34456
rect 27856 34416 27862 34428
rect 28445 34425 28457 34428
rect 28491 34425 28503 34459
rect 29638 34456 29644 34468
rect 29599 34428 29644 34456
rect 28445 34419 28503 34425
rect 29638 34416 29644 34428
rect 29696 34416 29702 34468
rect 18598 34388 18604 34400
rect 16908 34360 18604 34388
rect 16908 34348 16914 34360
rect 18598 34348 18604 34360
rect 18656 34348 18662 34400
rect 18693 34391 18751 34397
rect 18693 34357 18705 34391
rect 18739 34388 18751 34391
rect 19242 34388 19248 34400
rect 18739 34360 19248 34388
rect 18739 34357 18751 34360
rect 18693 34351 18751 34357
rect 19242 34348 19248 34360
rect 19300 34348 19306 34400
rect 19889 34391 19947 34397
rect 19889 34357 19901 34391
rect 19935 34388 19947 34391
rect 20438 34388 20444 34400
rect 19935 34360 20444 34388
rect 19935 34357 19947 34360
rect 19889 34351 19947 34357
rect 20438 34348 20444 34360
rect 20496 34348 20502 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 9398 34184 9404 34196
rect 9359 34156 9404 34184
rect 9398 34144 9404 34156
rect 9456 34144 9462 34196
rect 10686 34144 10692 34196
rect 10744 34184 10750 34196
rect 14458 34184 14464 34196
rect 10744 34156 14464 34184
rect 10744 34144 10750 34156
rect 14458 34144 14464 34156
rect 14516 34144 14522 34196
rect 15470 34144 15476 34196
rect 15528 34184 15534 34196
rect 16853 34187 16911 34193
rect 16853 34184 16865 34187
rect 15528 34156 16865 34184
rect 15528 34144 15534 34156
rect 16853 34153 16865 34156
rect 16899 34153 16911 34187
rect 16853 34147 16911 34153
rect 19426 34144 19432 34196
rect 19484 34184 19490 34196
rect 20530 34184 20536 34196
rect 19484 34156 20536 34184
rect 19484 34144 19490 34156
rect 20530 34144 20536 34156
rect 20588 34144 20594 34196
rect 23661 34187 23719 34193
rect 23661 34153 23673 34187
rect 23707 34184 23719 34187
rect 23842 34184 23848 34196
rect 23707 34156 23848 34184
rect 23707 34153 23719 34156
rect 23661 34147 23719 34153
rect 23842 34144 23848 34156
rect 23900 34144 23906 34196
rect 30561 34187 30619 34193
rect 30561 34153 30573 34187
rect 30607 34184 30619 34187
rect 30742 34184 30748 34196
rect 30607 34156 30748 34184
rect 30607 34153 30619 34156
rect 30561 34147 30619 34153
rect 30742 34144 30748 34156
rect 30800 34144 30806 34196
rect 31202 34184 31208 34196
rect 31163 34156 31208 34184
rect 31202 34144 31208 34156
rect 31260 34144 31266 34196
rect 9858 34076 9864 34128
rect 9916 34076 9922 34128
rect 10962 34076 10968 34128
rect 11020 34116 11026 34128
rect 13357 34119 13415 34125
rect 13357 34116 13369 34119
rect 11020 34088 13369 34116
rect 11020 34076 11026 34088
rect 13357 34085 13369 34088
rect 13403 34085 13415 34119
rect 16666 34116 16672 34128
rect 13357 34079 13415 34085
rect 16224 34088 16672 34116
rect 9876 34048 9904 34076
rect 10781 34051 10839 34057
rect 10781 34048 10793 34051
rect 9784 34020 10793 34048
rect 9784 33989 9812 34020
rect 10781 34017 10793 34020
rect 10827 34017 10839 34051
rect 14458 34048 14464 34060
rect 10781 34011 10839 34017
rect 12452 34020 14464 34048
rect 9677 33983 9735 33989
rect 9677 33949 9689 33983
rect 9723 33949 9735 33983
rect 9677 33943 9735 33949
rect 9769 33983 9827 33989
rect 9769 33949 9781 33983
rect 9815 33949 9827 33983
rect 9769 33943 9827 33949
rect 9861 33983 9919 33989
rect 9861 33949 9873 33983
rect 9907 33980 9919 33983
rect 9950 33980 9956 33992
rect 9907 33952 9956 33980
rect 9907 33949 9919 33952
rect 9861 33943 9919 33949
rect 9692 33912 9720 33943
rect 9950 33940 9956 33952
rect 10008 33940 10014 33992
rect 10045 33983 10103 33989
rect 10045 33949 10057 33983
rect 10091 33980 10103 33983
rect 10226 33980 10232 33992
rect 10091 33952 10232 33980
rect 10091 33949 10103 33952
rect 10045 33943 10103 33949
rect 10226 33940 10232 33952
rect 10284 33940 10290 33992
rect 10505 33983 10563 33989
rect 10505 33949 10517 33983
rect 10551 33980 10563 33983
rect 10686 33980 10692 33992
rect 10551 33952 10692 33980
rect 10551 33949 10563 33952
rect 10505 33943 10563 33949
rect 10686 33940 10692 33952
rect 10744 33940 10750 33992
rect 11974 33940 11980 33992
rect 12032 33980 12038 33992
rect 12342 33989 12348 33992
rect 12161 33983 12219 33989
rect 12161 33980 12173 33983
rect 12032 33952 12173 33980
rect 12032 33940 12038 33952
rect 12161 33949 12173 33952
rect 12207 33949 12219 33983
rect 12161 33943 12219 33949
rect 12309 33983 12348 33989
rect 12309 33949 12321 33983
rect 12309 33943 12348 33949
rect 12342 33940 12348 33943
rect 12400 33940 12406 33992
rect 12452 33989 12480 34020
rect 14458 34008 14464 34020
rect 14516 34048 14522 34060
rect 14516 34020 15240 34048
rect 14516 34008 14522 34020
rect 12437 33983 12495 33989
rect 12437 33949 12449 33983
rect 12483 33949 12495 33983
rect 12618 33980 12624 33992
rect 12577 33952 12624 33980
rect 12437 33943 12495 33949
rect 12618 33940 12624 33952
rect 12676 33989 12682 33992
rect 12676 33983 12725 33989
rect 12676 33949 12679 33983
rect 12713 33980 12725 33983
rect 12713 33952 13324 33980
rect 12713 33949 12725 33952
rect 12676 33943 12725 33949
rect 12676 33940 12682 33943
rect 11514 33912 11520 33924
rect 9692 33884 11520 33912
rect 11514 33872 11520 33884
rect 11572 33872 11578 33924
rect 12529 33915 12587 33921
rect 12529 33881 12541 33915
rect 12575 33912 12587 33915
rect 13078 33912 13084 33924
rect 12575 33884 13084 33912
rect 12575 33881 12587 33884
rect 12529 33875 12587 33881
rect 13078 33872 13084 33884
rect 13136 33872 13142 33924
rect 13296 33912 13324 33952
rect 13354 33940 13360 33992
rect 13412 33980 13418 33992
rect 15212 33989 15240 34020
rect 16224 33989 16252 34088
rect 16666 34076 16672 34088
rect 16724 34076 16730 34128
rect 18230 34076 18236 34128
rect 18288 34116 18294 34128
rect 29549 34119 29607 34125
rect 18288 34088 20990 34116
rect 18288 34076 18294 34088
rect 16758 34048 16764 34060
rect 16592 34020 16764 34048
rect 13541 33983 13599 33989
rect 13541 33980 13553 33983
rect 13412 33952 13553 33980
rect 13412 33940 13418 33952
rect 13541 33949 13553 33952
rect 13587 33949 13599 33983
rect 13541 33943 13599 33949
rect 14921 33983 14979 33989
rect 14921 33949 14933 33983
rect 14967 33949 14979 33983
rect 14921 33943 14979 33949
rect 15197 33983 15255 33989
rect 15197 33949 15209 33983
rect 15243 33949 15255 33983
rect 15197 33943 15255 33949
rect 16209 33983 16267 33989
rect 16209 33949 16221 33983
rect 16255 33949 16267 33983
rect 16209 33943 16267 33949
rect 16302 33983 16360 33989
rect 16302 33949 16314 33983
rect 16348 33949 16360 33983
rect 16482 33980 16488 33992
rect 16443 33952 16488 33980
rect 16302 33943 16360 33949
rect 14936 33912 14964 33943
rect 15562 33912 15568 33924
rect 13296 33884 14403 33912
rect 14936 33884 15568 33912
rect 12618 33804 12624 33856
rect 12676 33844 12682 33856
rect 12805 33847 12863 33853
rect 12805 33844 12817 33847
rect 12676 33816 12817 33844
rect 12676 33804 12682 33816
rect 12805 33813 12817 33816
rect 12851 33813 12863 33847
rect 12805 33807 12863 33813
rect 13814 33804 13820 33856
rect 13872 33844 13878 33856
rect 14274 33844 14280 33856
rect 13872 33816 14280 33844
rect 13872 33804 13878 33816
rect 14274 33804 14280 33816
rect 14332 33804 14338 33856
rect 14375 33844 14403 33884
rect 15562 33872 15568 33884
rect 15620 33872 15626 33924
rect 16316 33912 16344 33943
rect 16482 33940 16488 33952
rect 16540 33940 16546 33992
rect 16592 33989 16620 34020
rect 16758 34008 16764 34020
rect 16816 34008 16822 34060
rect 16577 33983 16635 33989
rect 16577 33949 16589 33983
rect 16623 33949 16635 33983
rect 16577 33943 16635 33949
rect 16666 33940 16672 33992
rect 16724 33989 16730 33992
rect 16724 33980 16732 33989
rect 17402 33980 17408 33992
rect 16724 33952 16769 33980
rect 17363 33952 17408 33980
rect 16724 33943 16732 33952
rect 16724 33940 16730 33943
rect 17402 33940 17408 33952
rect 17460 33940 17466 33992
rect 17681 33983 17739 33989
rect 17681 33949 17693 33983
rect 17727 33980 17739 33983
rect 17954 33980 17960 33992
rect 17727 33952 17960 33980
rect 17727 33949 17739 33952
rect 17681 33943 17739 33949
rect 17954 33940 17960 33952
rect 18012 33940 18018 33992
rect 19242 33980 19248 33992
rect 19203 33952 19248 33980
rect 19242 33940 19248 33952
rect 19300 33940 19306 33992
rect 19426 33989 19432 33992
rect 19393 33983 19432 33989
rect 19393 33949 19405 33983
rect 19393 33943 19432 33949
rect 19426 33940 19432 33943
rect 19484 33940 19490 33992
rect 19749 33983 19807 33989
rect 19749 33949 19761 33983
rect 19795 33980 19807 33983
rect 19904 33980 19932 34088
rect 20070 34008 20076 34060
rect 20128 34008 20134 34060
rect 20714 34008 20720 34060
rect 20772 34008 20778 34060
rect 20962 34048 20990 34088
rect 29549 34085 29561 34119
rect 29595 34116 29607 34119
rect 30190 34116 30196 34128
rect 29595 34088 30196 34116
rect 29595 34085 29607 34088
rect 29549 34079 29607 34085
rect 30190 34076 30196 34088
rect 30248 34076 30254 34128
rect 20962 34020 22145 34048
rect 19795 33952 19932 33980
rect 19795 33949 19807 33952
rect 19749 33943 19807 33949
rect 16942 33912 16948 33924
rect 16316 33884 16948 33912
rect 16942 33872 16948 33884
rect 17000 33872 17006 33924
rect 17862 33872 17868 33924
rect 17920 33912 17926 33924
rect 19058 33912 19064 33924
rect 17920 33884 19064 33912
rect 17920 33872 17926 33884
rect 19058 33872 19064 33884
rect 19116 33912 19122 33924
rect 19521 33915 19579 33921
rect 19521 33912 19533 33915
rect 19116 33884 19533 33912
rect 19116 33872 19122 33884
rect 19521 33881 19533 33884
rect 19567 33881 19579 33915
rect 19521 33875 19579 33881
rect 19618 33872 19624 33924
rect 19676 33921 19682 33924
rect 19676 33915 19691 33921
rect 19679 33881 19691 33915
rect 20088 33912 20116 34008
rect 20438 33980 20444 33992
rect 20399 33952 20444 33980
rect 20438 33940 20444 33952
rect 20496 33940 20502 33992
rect 20530 33940 20536 33992
rect 20588 33980 20594 33992
rect 20732 33980 20760 34008
rect 20962 33989 20990 34020
rect 20809 33983 20867 33989
rect 20809 33980 20821 33983
rect 20588 33952 20633 33980
rect 20732 33952 20821 33980
rect 20588 33940 20594 33952
rect 20809 33949 20821 33952
rect 20855 33949 20867 33983
rect 20809 33943 20867 33949
rect 20947 33983 21005 33989
rect 20947 33949 20959 33983
rect 20993 33949 21005 33983
rect 21634 33980 21640 33992
rect 21595 33952 21640 33980
rect 20947 33943 21005 33949
rect 21634 33940 21640 33952
rect 21692 33940 21698 33992
rect 21818 33989 21824 33992
rect 21785 33983 21824 33989
rect 21785 33949 21797 33983
rect 21785 33943 21824 33949
rect 21818 33940 21824 33943
rect 21876 33940 21882 33992
rect 22002 33980 22008 33992
rect 21963 33952 22008 33980
rect 22002 33940 22008 33952
rect 22060 33940 22066 33992
rect 22117 33989 22145 34020
rect 22102 33983 22160 33989
rect 22102 33949 22114 33983
rect 22148 33949 22160 33983
rect 23290 33980 23296 33992
rect 23251 33952 23296 33980
rect 22102 33943 22160 33949
rect 23290 33940 23296 33952
rect 23348 33940 23354 33992
rect 24581 33983 24639 33989
rect 24581 33980 24593 33983
rect 23860 33952 24593 33980
rect 20717 33915 20775 33921
rect 20717 33912 20729 33915
rect 20088 33884 20729 33912
rect 19676 33875 19691 33881
rect 20717 33881 20729 33884
rect 20763 33912 20775 33915
rect 21913 33915 21971 33921
rect 21913 33912 21925 33915
rect 20763 33884 21925 33912
rect 20763 33881 20775 33884
rect 20717 33875 20775 33881
rect 21913 33881 21925 33884
rect 21959 33881 21971 33915
rect 21913 33875 21971 33881
rect 19676 33872 19682 33875
rect 15102 33844 15108 33856
rect 14375 33816 15108 33844
rect 15102 33804 15108 33816
rect 15160 33804 15166 33856
rect 16666 33804 16672 33856
rect 16724 33844 16730 33856
rect 17310 33844 17316 33856
rect 16724 33816 17316 33844
rect 16724 33804 16730 33816
rect 17310 33804 17316 33816
rect 17368 33844 17374 33856
rect 18230 33844 18236 33856
rect 17368 33816 18236 33844
rect 17368 33804 17374 33816
rect 18230 33804 18236 33816
rect 18288 33804 18294 33856
rect 19889 33847 19947 33853
rect 19889 33813 19901 33847
rect 19935 33844 19947 33847
rect 19978 33844 19984 33856
rect 19935 33816 19984 33844
rect 19935 33813 19947 33816
rect 19889 33807 19947 33813
rect 19978 33804 19984 33816
rect 20036 33804 20042 33856
rect 21082 33844 21088 33856
rect 21043 33816 21088 33844
rect 21082 33804 21088 33816
rect 21140 33804 21146 33856
rect 22281 33847 22339 33853
rect 22281 33813 22293 33847
rect 22327 33844 22339 33847
rect 22462 33844 22468 33856
rect 22327 33816 22468 33844
rect 22327 33813 22339 33816
rect 22281 33807 22339 33813
rect 22462 33804 22468 33816
rect 22520 33804 22526 33856
rect 23658 33844 23664 33856
rect 23619 33816 23664 33844
rect 23658 33804 23664 33816
rect 23716 33804 23722 33856
rect 23860 33853 23888 33952
rect 24581 33949 24593 33952
rect 24627 33949 24639 33983
rect 28074 33980 28080 33992
rect 28035 33952 28080 33980
rect 24581 33943 24639 33949
rect 28074 33940 28080 33952
rect 28132 33940 28138 33992
rect 29546 33980 29552 33992
rect 29507 33952 29552 33980
rect 29546 33940 29552 33952
rect 29604 33940 29610 33992
rect 29733 33983 29791 33989
rect 29733 33949 29745 33983
rect 29779 33980 29791 33983
rect 30558 33980 30564 33992
rect 29779 33952 30564 33980
rect 29779 33949 29791 33952
rect 29733 33943 29791 33949
rect 30558 33940 30564 33952
rect 30616 33940 30622 33992
rect 31389 33983 31447 33989
rect 31389 33980 31401 33983
rect 30760 33952 31401 33980
rect 24762 33872 24768 33924
rect 24820 33912 24826 33924
rect 25685 33915 25743 33921
rect 25685 33912 25697 33915
rect 24820 33884 25697 33912
rect 24820 33872 24826 33884
rect 25685 33881 25697 33884
rect 25731 33912 25743 33915
rect 26510 33912 26516 33924
rect 25731 33884 26516 33912
rect 25731 33881 25743 33884
rect 25685 33875 25743 33881
rect 26510 33872 26516 33884
rect 26568 33872 26574 33924
rect 23845 33847 23903 33853
rect 23845 33813 23857 33847
rect 23891 33813 23903 33847
rect 23845 33807 23903 33813
rect 24026 33804 24032 33856
rect 24084 33844 24090 33856
rect 24397 33847 24455 33853
rect 24397 33844 24409 33847
rect 24084 33816 24409 33844
rect 24084 33804 24090 33816
rect 24397 33813 24409 33816
rect 24443 33813 24455 33847
rect 24397 33807 24455 33813
rect 25038 33804 25044 33856
rect 25096 33844 25102 33856
rect 26973 33847 27031 33853
rect 26973 33844 26985 33847
rect 25096 33816 26985 33844
rect 25096 33804 25102 33816
rect 26973 33813 26985 33816
rect 27019 33844 27031 33847
rect 27522 33844 27528 33856
rect 27019 33816 27528 33844
rect 27019 33813 27031 33816
rect 26973 33807 27031 33813
rect 27522 33804 27528 33816
rect 27580 33804 27586 33856
rect 27890 33844 27896 33856
rect 27851 33816 27896 33844
rect 27890 33804 27896 33816
rect 27948 33804 27954 33856
rect 30282 33804 30288 33856
rect 30340 33844 30346 33856
rect 30760 33853 30788 33952
rect 31389 33949 31401 33952
rect 31435 33949 31447 33983
rect 31389 33943 31447 33949
rect 30561 33847 30619 33853
rect 30561 33844 30573 33847
rect 30340 33816 30573 33844
rect 30340 33804 30346 33816
rect 30561 33813 30573 33816
rect 30607 33813 30619 33847
rect 30561 33807 30619 33813
rect 30745 33847 30803 33853
rect 30745 33813 30757 33847
rect 30791 33813 30803 33847
rect 30745 33807 30803 33813
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 10410 33640 10416 33652
rect 10371 33612 10416 33640
rect 10410 33600 10416 33612
rect 10468 33600 10474 33652
rect 11974 33640 11980 33652
rect 11935 33612 11980 33640
rect 11974 33600 11980 33612
rect 12032 33600 12038 33652
rect 12158 33600 12164 33652
rect 12216 33640 12222 33652
rect 13630 33640 13636 33652
rect 12216 33612 12388 33640
rect 13591 33612 13636 33640
rect 12216 33600 12222 33612
rect 10045 33575 10103 33581
rect 10045 33541 10057 33575
rect 10091 33572 10103 33575
rect 10778 33572 10784 33584
rect 10091 33544 10784 33572
rect 10091 33541 10103 33544
rect 10045 33535 10103 33541
rect 10778 33532 10784 33544
rect 10836 33572 10842 33584
rect 10962 33572 10968 33584
rect 10836 33544 10968 33572
rect 10836 33532 10842 33544
rect 10962 33532 10968 33544
rect 11020 33532 11026 33584
rect 11054 33532 11060 33584
rect 11112 33572 11118 33584
rect 12360 33581 12388 33612
rect 13630 33600 13636 33612
rect 13688 33600 13694 33652
rect 15933 33643 15991 33649
rect 15933 33640 15945 33643
rect 13740 33612 15945 33640
rect 12345 33575 12403 33581
rect 12345 33572 12357 33575
rect 11112 33544 12357 33572
rect 11112 33532 11118 33544
rect 12345 33541 12357 33544
rect 12391 33541 12403 33575
rect 12345 33535 12403 33541
rect 12434 33532 12440 33584
rect 12492 33581 12498 33584
rect 12492 33575 12521 33581
rect 12509 33541 12521 33575
rect 12492 33535 12521 33541
rect 12492 33532 12498 33535
rect 13538 33532 13544 33584
rect 13596 33572 13602 33584
rect 13740 33572 13768 33612
rect 15933 33609 15945 33612
rect 15979 33609 15991 33643
rect 15933 33603 15991 33609
rect 16482 33600 16488 33652
rect 16540 33640 16546 33652
rect 17862 33640 17868 33652
rect 16540 33612 17868 33640
rect 16540 33600 16546 33612
rect 17862 33600 17868 33612
rect 17920 33600 17926 33652
rect 18322 33600 18328 33652
rect 18380 33640 18386 33652
rect 18690 33640 18696 33652
rect 18380 33612 18696 33640
rect 18380 33600 18386 33612
rect 18690 33600 18696 33612
rect 18748 33640 18754 33652
rect 20438 33640 20444 33652
rect 18748 33612 20444 33640
rect 18748 33600 18754 33612
rect 20438 33600 20444 33612
rect 20496 33600 20502 33652
rect 20533 33643 20591 33649
rect 20533 33609 20545 33643
rect 20579 33640 20591 33643
rect 21634 33640 21640 33652
rect 20579 33612 21640 33640
rect 20579 33609 20591 33612
rect 20533 33603 20591 33609
rect 21634 33600 21640 33612
rect 21692 33600 21698 33652
rect 23290 33600 23296 33652
rect 23348 33640 23354 33652
rect 24213 33643 24271 33649
rect 24213 33640 24225 33643
rect 23348 33612 24225 33640
rect 23348 33600 23354 33612
rect 24213 33609 24225 33612
rect 24259 33609 24271 33643
rect 26421 33643 26479 33649
rect 26421 33640 26433 33643
rect 24213 33603 24271 33609
rect 24320 33612 26433 33640
rect 13596 33544 13768 33572
rect 14139 33575 14197 33581
rect 13596 33532 13602 33544
rect 14139 33541 14151 33575
rect 14185 33572 14197 33575
rect 14274 33572 14280 33584
rect 14185 33544 14280 33572
rect 14185 33541 14197 33544
rect 14139 33535 14197 33541
rect 14274 33532 14280 33544
rect 14332 33532 14338 33584
rect 14826 33572 14832 33584
rect 14384 33544 14832 33572
rect 10229 33507 10287 33513
rect 10229 33473 10241 33507
rect 10275 33504 10287 33507
rect 10594 33504 10600 33516
rect 10275 33476 10600 33504
rect 10275 33473 10287 33476
rect 10229 33467 10287 33473
rect 10594 33464 10600 33476
rect 10652 33464 10658 33516
rect 12158 33504 12164 33516
rect 12119 33476 12164 33504
rect 12158 33464 12164 33476
rect 12216 33464 12222 33516
rect 12253 33507 12311 33513
rect 12253 33473 12265 33507
rect 12299 33473 12311 33507
rect 12253 33467 12311 33473
rect 12268 33436 12296 33467
rect 13630 33464 13636 33516
rect 13688 33510 13694 33516
rect 13817 33510 13875 33513
rect 13688 33507 13875 33510
rect 13688 33482 13829 33507
rect 13688 33464 13694 33482
rect 13796 33476 13829 33482
rect 13817 33473 13829 33476
rect 13863 33473 13875 33507
rect 13817 33467 13875 33473
rect 13909 33507 13967 33513
rect 13909 33473 13921 33507
rect 13955 33473 13967 33507
rect 13909 33467 13967 33473
rect 14001 33507 14059 33513
rect 14001 33473 14013 33507
rect 14047 33504 14059 33507
rect 14384 33504 14412 33544
rect 14826 33532 14832 33544
rect 14884 33532 14890 33584
rect 15378 33572 15384 33584
rect 14936 33544 15384 33572
rect 14936 33516 14964 33544
rect 15378 33532 15384 33544
rect 15436 33532 15442 33584
rect 16942 33532 16948 33584
rect 17000 33572 17006 33584
rect 17126 33572 17132 33584
rect 17000 33544 17132 33572
rect 17000 33532 17006 33544
rect 17126 33532 17132 33544
rect 17184 33532 17190 33584
rect 18966 33532 18972 33584
rect 19024 33572 19030 33584
rect 20809 33575 20867 33581
rect 20809 33572 20821 33575
rect 19024 33544 20821 33572
rect 19024 33532 19030 33544
rect 20809 33541 20821 33544
rect 20855 33541 20867 33575
rect 20809 33535 20867 33541
rect 20901 33575 20959 33581
rect 20901 33541 20913 33575
rect 20947 33572 20959 33575
rect 21542 33572 21548 33584
rect 20947 33544 21548 33572
rect 20947 33541 20959 33544
rect 20901 33535 20959 33541
rect 21542 33532 21548 33544
rect 21600 33532 21606 33584
rect 21818 33532 21824 33584
rect 21876 33572 21882 33584
rect 24320 33572 24348 33612
rect 26421 33609 26433 33612
rect 26467 33609 26479 33643
rect 26421 33603 26479 33609
rect 26510 33600 26516 33652
rect 26568 33640 26574 33652
rect 27246 33640 27252 33652
rect 26568 33612 27252 33640
rect 26568 33600 26574 33612
rect 27246 33600 27252 33612
rect 27304 33640 27310 33652
rect 29549 33643 29607 33649
rect 29549 33640 29561 33643
rect 27304 33612 29561 33640
rect 27304 33600 27310 33612
rect 29549 33609 29561 33612
rect 29595 33640 29607 33643
rect 30374 33640 30380 33652
rect 29595 33612 30380 33640
rect 29595 33609 29607 33612
rect 29549 33603 29607 33609
rect 30374 33600 30380 33612
rect 30432 33600 30438 33652
rect 21876 33544 24348 33572
rect 25308 33575 25366 33581
rect 21876 33532 21882 33544
rect 25308 33541 25320 33575
rect 25354 33572 25366 33575
rect 27890 33572 27896 33584
rect 25354 33544 27896 33572
rect 25354 33541 25366 33544
rect 25308 33535 25366 33541
rect 27890 33532 27896 33544
rect 27948 33532 27954 33584
rect 30282 33572 30288 33584
rect 30243 33544 30288 33572
rect 30282 33532 30288 33544
rect 30340 33532 30346 33584
rect 14918 33504 14924 33516
rect 14047 33476 14412 33504
rect 14831 33476 14924 33504
rect 14047 33473 14059 33476
rect 14001 33467 14059 33473
rect 12342 33436 12348 33448
rect 12268 33408 12348 33436
rect 12342 33396 12348 33408
rect 12400 33396 12406 33448
rect 12621 33439 12679 33445
rect 12621 33405 12633 33439
rect 12667 33436 12679 33439
rect 12710 33436 12716 33448
rect 12667 33408 12716 33436
rect 12667 33405 12679 33408
rect 12621 33399 12679 33405
rect 12710 33396 12716 33408
rect 12768 33396 12774 33448
rect 13924 33436 13952 33467
rect 14918 33464 14924 33476
rect 14976 33464 14982 33516
rect 15013 33507 15071 33513
rect 15013 33473 15025 33507
rect 15059 33473 15071 33507
rect 15013 33467 15071 33473
rect 15105 33507 15163 33513
rect 15105 33473 15117 33507
rect 15151 33473 15163 33507
rect 15105 33467 15163 33473
rect 15243 33507 15301 33513
rect 15243 33473 15255 33507
rect 15289 33504 15301 33507
rect 15838 33504 15844 33516
rect 15289 33476 15844 33504
rect 15289 33473 15301 33476
rect 15243 33467 15301 33473
rect 14277 33439 14335 33445
rect 13924 33408 14044 33436
rect 14016 33368 14044 33408
rect 14277 33405 14289 33439
rect 14323 33436 14335 33439
rect 14826 33436 14832 33448
rect 14323 33408 14832 33436
rect 14323 33405 14335 33408
rect 14277 33399 14335 33405
rect 14826 33396 14832 33408
rect 14884 33396 14890 33448
rect 15028 33436 15056 33467
rect 14936 33408 15056 33436
rect 14936 33380 14964 33408
rect 14016 33340 14320 33368
rect 14292 33312 14320 33340
rect 14918 33328 14924 33380
rect 14976 33328 14982 33380
rect 15010 33328 15016 33380
rect 15068 33368 15074 33380
rect 15120 33368 15148 33467
rect 15838 33464 15844 33476
rect 15896 33464 15902 33516
rect 16025 33507 16083 33513
rect 16025 33473 16037 33507
rect 16071 33504 16083 33507
rect 18138 33504 18144 33516
rect 16071 33476 18144 33504
rect 16071 33473 16083 33476
rect 16025 33467 16083 33473
rect 18138 33464 18144 33476
rect 18196 33464 18202 33516
rect 18230 33464 18236 33516
rect 18288 33504 18294 33516
rect 18288 33476 18333 33504
rect 18288 33464 18294 33476
rect 18598 33464 18604 33516
rect 18656 33504 18662 33516
rect 20717 33507 20775 33513
rect 20717 33504 20729 33507
rect 18656 33476 20729 33504
rect 18656 33464 18662 33476
rect 20717 33473 20729 33476
rect 20763 33473 20775 33507
rect 20717 33467 20775 33473
rect 20990 33464 20996 33516
rect 21048 33513 21054 33516
rect 21048 33507 21077 33513
rect 21065 33473 21077 33507
rect 21048 33467 21077 33473
rect 21048 33464 21054 33467
rect 22278 33464 22284 33516
rect 22336 33504 22342 33516
rect 22445 33507 22503 33513
rect 22445 33504 22457 33507
rect 22336 33476 22457 33504
rect 22336 33464 22342 33476
rect 22445 33473 22457 33476
rect 22491 33473 22503 33507
rect 24118 33504 24124 33516
rect 24079 33476 24124 33504
rect 22445 33467 22503 33473
rect 24118 33464 24124 33476
rect 24176 33464 24182 33516
rect 24305 33507 24363 33513
rect 24305 33473 24317 33507
rect 24351 33504 24363 33507
rect 24578 33504 24584 33516
rect 24351 33476 24584 33504
rect 24351 33473 24363 33476
rect 24305 33467 24363 33473
rect 24578 33464 24584 33476
rect 24636 33464 24642 33516
rect 25038 33504 25044 33516
rect 24999 33476 25044 33504
rect 25038 33464 25044 33476
rect 25096 33464 25102 33516
rect 27522 33504 27528 33516
rect 27483 33476 27528 33504
rect 27522 33464 27528 33476
rect 27580 33464 27586 33516
rect 27798 33513 27804 33516
rect 27792 33467 27804 33513
rect 27856 33504 27862 33516
rect 27856 33476 27892 33504
rect 27798 33464 27804 33467
rect 27856 33464 27862 33476
rect 28994 33464 29000 33516
rect 29052 33504 29058 33516
rect 29457 33507 29515 33513
rect 29457 33504 29469 33507
rect 29052 33476 29469 33504
rect 29052 33464 29058 33476
rect 29457 33473 29469 33476
rect 29503 33473 29515 33507
rect 29457 33467 29515 33473
rect 29546 33464 29552 33516
rect 29604 33504 29610 33516
rect 30193 33507 30251 33513
rect 30193 33504 30205 33507
rect 29604 33476 30205 33504
rect 29604 33464 29610 33476
rect 30193 33473 30205 33476
rect 30239 33473 30251 33507
rect 30193 33467 30251 33473
rect 30377 33507 30435 33513
rect 30377 33473 30389 33507
rect 30423 33504 30435 33507
rect 30558 33504 30564 33516
rect 30423 33476 30564 33504
rect 30423 33473 30435 33476
rect 30377 33467 30435 33473
rect 30558 33464 30564 33476
rect 30616 33504 30622 33516
rect 30834 33504 30840 33516
rect 30616 33476 30840 33504
rect 30616 33464 30622 33476
rect 30834 33464 30840 33476
rect 30892 33464 30898 33516
rect 15381 33439 15439 33445
rect 15381 33405 15393 33439
rect 15427 33436 15439 33439
rect 16206 33436 16212 33448
rect 15427 33408 16212 33436
rect 15427 33405 15439 33408
rect 15381 33399 15439 33405
rect 15068 33340 15148 33368
rect 15068 33328 15074 33340
rect 14274 33260 14280 33312
rect 14332 33260 14338 33312
rect 14642 33260 14648 33312
rect 14700 33300 14706 33312
rect 14737 33303 14795 33309
rect 14737 33300 14749 33303
rect 14700 33272 14749 33300
rect 14700 33260 14706 33272
rect 14737 33269 14749 33272
rect 14783 33269 14795 33303
rect 14737 33263 14795 33269
rect 14826 33260 14832 33312
rect 14884 33300 14890 33312
rect 15396 33300 15424 33399
rect 16206 33396 16212 33408
rect 16264 33396 16270 33448
rect 16666 33436 16672 33448
rect 16627 33408 16672 33436
rect 16666 33396 16672 33408
rect 16724 33396 16730 33448
rect 16850 33396 16856 33448
rect 16908 33436 16914 33448
rect 16945 33439 17003 33445
rect 16945 33436 16957 33439
rect 16908 33408 16957 33436
rect 16908 33396 16914 33408
rect 16945 33405 16957 33408
rect 16991 33405 17003 33439
rect 16945 33399 17003 33405
rect 17770 33396 17776 33448
rect 17828 33436 17834 33448
rect 17957 33439 18015 33445
rect 17957 33436 17969 33439
rect 17828 33408 17969 33436
rect 17828 33396 17834 33408
rect 17957 33405 17969 33408
rect 18003 33405 18015 33439
rect 17957 33399 18015 33405
rect 18046 33396 18052 33448
rect 18104 33436 18110 33448
rect 18616 33436 18644 33464
rect 18104 33408 18644 33436
rect 19245 33439 19303 33445
rect 18104 33396 18110 33408
rect 19245 33405 19257 33439
rect 19291 33436 19303 33439
rect 20346 33436 20352 33448
rect 19291 33408 20352 33436
rect 19291 33405 19303 33408
rect 19245 33399 19303 33405
rect 20346 33396 20352 33408
rect 20404 33396 20410 33448
rect 20438 33396 20444 33448
rect 20496 33396 20502 33448
rect 20898 33396 20904 33448
rect 20956 33436 20962 33448
rect 21177 33439 21235 33445
rect 21177 33436 21189 33439
rect 20956 33408 21189 33436
rect 20956 33396 20962 33408
rect 21177 33405 21189 33408
rect 21223 33405 21235 33439
rect 22186 33436 22192 33448
rect 22147 33408 22192 33436
rect 21177 33399 21235 33405
rect 22186 33396 22192 33408
rect 22244 33396 22250 33448
rect 19475 33371 19533 33377
rect 19475 33337 19487 33371
rect 19521 33368 19533 33371
rect 20456 33368 20484 33396
rect 20916 33368 20944 33396
rect 19521 33340 20944 33368
rect 19521 33337 19533 33340
rect 19475 33331 19533 33337
rect 14884 33272 15424 33300
rect 14884 33260 14890 33272
rect 23474 33260 23480 33312
rect 23532 33300 23538 33312
rect 23569 33303 23627 33309
rect 23569 33300 23581 33303
rect 23532 33272 23581 33300
rect 23532 33260 23538 33272
rect 23569 33269 23581 33272
rect 23615 33269 23627 33303
rect 23569 33263 23627 33269
rect 28534 33260 28540 33312
rect 28592 33300 28598 33312
rect 28905 33303 28963 33309
rect 28905 33300 28917 33303
rect 28592 33272 28917 33300
rect 28592 33260 28598 33272
rect 28905 33269 28917 33272
rect 28951 33269 28963 33303
rect 28905 33263 28963 33269
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 18322 33096 18328 33108
rect 9048 33068 18328 33096
rect 9048 32901 9076 33068
rect 18322 33056 18328 33068
rect 18380 33056 18386 33108
rect 19334 33056 19340 33108
rect 19392 33096 19398 33108
rect 20070 33096 20076 33108
rect 19392 33068 20076 33096
rect 19392 33056 19398 33068
rect 20070 33056 20076 33068
rect 20128 33056 20134 33108
rect 21913 33099 21971 33105
rect 21913 33065 21925 33099
rect 21959 33096 21971 33099
rect 22278 33096 22284 33108
rect 21959 33068 22284 33096
rect 21959 33065 21971 33068
rect 21913 33059 21971 33065
rect 22278 33056 22284 33068
rect 22336 33056 22342 33108
rect 28718 33056 28724 33108
rect 28776 33096 28782 33108
rect 28997 33099 29055 33105
rect 28997 33096 29009 33099
rect 28776 33068 29009 33096
rect 28776 33056 28782 33068
rect 28997 33065 29009 33068
rect 29043 33065 29055 33099
rect 28997 33059 29055 33065
rect 9950 32988 9956 33040
rect 10008 32988 10014 33040
rect 12066 33028 12072 33040
rect 12027 33000 12072 33028
rect 12066 32988 12072 33000
rect 12124 32988 12130 33040
rect 13262 32988 13268 33040
rect 13320 33028 13326 33040
rect 13320 33000 14136 33028
rect 13320 32988 13326 33000
rect 9968 32960 9996 32988
rect 11149 32963 11207 32969
rect 11149 32960 11161 32963
rect 9968 32932 10088 32960
rect 10060 32901 10088 32932
rect 10152 32932 11161 32960
rect 10152 32901 10180 32932
rect 11149 32929 11161 32932
rect 11195 32929 11207 32963
rect 11149 32923 11207 32929
rect 12158 32920 12164 32972
rect 12216 32960 12222 32972
rect 13630 32960 13636 32972
rect 12216 32932 13636 32960
rect 12216 32920 12222 32932
rect 9033 32895 9091 32901
rect 9033 32861 9045 32895
rect 9079 32861 9091 32895
rect 9033 32855 9091 32861
rect 9953 32895 10011 32901
rect 9953 32861 9965 32895
rect 9999 32861 10011 32895
rect 9953 32855 10011 32861
rect 10042 32895 10100 32901
rect 10042 32861 10054 32895
rect 10088 32861 10100 32895
rect 10042 32855 10100 32861
rect 10137 32895 10195 32901
rect 10137 32861 10149 32895
rect 10183 32861 10195 32895
rect 10137 32855 10195 32861
rect 9217 32827 9275 32833
rect 9217 32793 9229 32827
rect 9263 32824 9275 32827
rect 9490 32824 9496 32836
rect 9263 32796 9496 32824
rect 9263 32793 9275 32796
rect 9217 32787 9275 32793
rect 9490 32784 9496 32796
rect 9548 32784 9554 32836
rect 9674 32756 9680 32768
rect 9635 32728 9680 32756
rect 9674 32716 9680 32728
rect 9732 32716 9738 32768
rect 9968 32756 9996 32855
rect 10226 32852 10232 32904
rect 10284 32892 10290 32904
rect 10321 32895 10379 32901
rect 10321 32892 10333 32895
rect 10284 32864 10333 32892
rect 10284 32852 10290 32864
rect 10321 32861 10333 32864
rect 10367 32861 10379 32895
rect 10778 32892 10784 32904
rect 10739 32864 10784 32892
rect 10321 32855 10379 32861
rect 10778 32852 10784 32864
rect 10836 32852 10842 32904
rect 10965 32895 11023 32901
rect 10965 32861 10977 32895
rect 11011 32892 11023 32895
rect 11054 32892 11060 32904
rect 11011 32864 11060 32892
rect 11011 32861 11023 32864
rect 10965 32855 11023 32861
rect 11054 32852 11060 32864
rect 11112 32852 11118 32904
rect 12268 32901 12296 32932
rect 13630 32920 13636 32932
rect 13688 32920 13694 32972
rect 14108 32969 14136 33000
rect 15562 32988 15568 33040
rect 15620 33028 15626 33040
rect 20441 33031 20499 33037
rect 15620 33000 17632 33028
rect 15620 32988 15626 33000
rect 14093 32963 14151 32969
rect 14093 32929 14105 32963
rect 14139 32929 14151 32963
rect 14093 32923 14151 32929
rect 16209 32963 16267 32969
rect 16209 32929 16221 32963
rect 16255 32960 16267 32963
rect 17402 32960 17408 32972
rect 16255 32932 17408 32960
rect 16255 32929 16267 32932
rect 16209 32923 16267 32929
rect 12253 32895 12311 32901
rect 12253 32861 12265 32895
rect 12299 32861 12311 32895
rect 12253 32855 12311 32861
rect 12342 32852 12348 32904
rect 12400 32892 12406 32904
rect 12710 32892 12716 32904
rect 12400 32864 12445 32892
rect 12623 32864 12716 32892
rect 12400 32852 12406 32864
rect 12710 32852 12716 32864
rect 12768 32892 12774 32904
rect 13354 32892 13360 32904
rect 12768 32864 13360 32892
rect 12768 32852 12774 32864
rect 13354 32852 13360 32864
rect 13412 32852 13418 32904
rect 14108 32892 14136 32923
rect 17402 32920 17408 32932
rect 17460 32920 17466 32972
rect 14182 32892 14188 32904
rect 14108 32864 14188 32892
rect 14182 32852 14188 32864
rect 14240 32852 14246 32904
rect 14918 32852 14924 32904
rect 14976 32892 14982 32904
rect 15654 32892 15660 32904
rect 14976 32864 15660 32892
rect 14976 32852 14982 32864
rect 15654 32852 15660 32864
rect 15712 32892 15718 32904
rect 17604 32901 17632 33000
rect 20441 32997 20453 33031
rect 20487 33028 20499 33031
rect 20530 33028 20536 33040
rect 20487 33000 20536 33028
rect 20487 32997 20499 33000
rect 20441 32991 20499 32997
rect 20530 32988 20536 33000
rect 20588 32988 20594 33040
rect 17862 32960 17868 32972
rect 17823 32932 17868 32960
rect 17862 32920 17868 32932
rect 17920 32920 17926 32972
rect 20180 32932 23612 32960
rect 16485 32895 16543 32901
rect 16485 32892 16497 32895
rect 15712 32864 16497 32892
rect 15712 32852 15718 32864
rect 16485 32861 16497 32864
rect 16531 32861 16543 32895
rect 16485 32855 16543 32861
rect 17589 32895 17647 32901
rect 17589 32861 17601 32895
rect 17635 32892 17647 32895
rect 18598 32892 18604 32904
rect 17635 32864 18604 32892
rect 17635 32861 17647 32864
rect 17589 32855 17647 32861
rect 18598 32852 18604 32864
rect 18656 32852 18662 32904
rect 19242 32892 19248 32904
rect 19203 32864 19248 32892
rect 19242 32852 19248 32864
rect 19300 32852 19306 32904
rect 19426 32892 19432 32904
rect 19387 32864 19432 32892
rect 19426 32852 19432 32864
rect 19484 32852 19490 32904
rect 19518 32852 19524 32904
rect 19576 32892 19582 32904
rect 19613 32895 19671 32901
rect 19613 32892 19625 32895
rect 19576 32864 19625 32892
rect 19576 32852 19582 32864
rect 19613 32861 19625 32864
rect 19659 32861 19671 32895
rect 19613 32855 19671 32861
rect 19702 32852 19708 32904
rect 19760 32892 19766 32904
rect 19760 32864 19805 32892
rect 19760 32852 19766 32864
rect 10594 32784 10600 32836
rect 10652 32824 10658 32836
rect 12437 32827 12495 32833
rect 10652 32796 12020 32824
rect 10652 32784 10658 32796
rect 11882 32756 11888 32768
rect 9968 32728 11888 32756
rect 11882 32716 11888 32728
rect 11940 32716 11946 32768
rect 11992 32756 12020 32796
rect 12437 32793 12449 32827
rect 12483 32793 12495 32827
rect 12437 32787 12495 32793
rect 12575 32827 12633 32833
rect 12575 32793 12587 32827
rect 12621 32824 12633 32827
rect 12802 32824 12808 32836
rect 12621 32796 12808 32824
rect 12621 32793 12633 32796
rect 12575 32787 12633 32793
rect 12452 32756 12480 32787
rect 12802 32784 12808 32796
rect 12860 32784 12866 32836
rect 14360 32827 14418 32833
rect 14360 32793 14372 32827
rect 14406 32824 14418 32827
rect 18230 32824 18236 32836
rect 14406 32796 18236 32824
rect 14406 32793 14418 32796
rect 14360 32787 14418 32793
rect 18230 32784 18236 32796
rect 18288 32784 18294 32836
rect 20180 32824 20208 32932
rect 22094 32892 22100 32904
rect 22055 32864 22100 32892
rect 22094 32852 22100 32864
rect 22152 32852 22158 32904
rect 22373 32895 22431 32901
rect 22373 32861 22385 32895
rect 22419 32892 22431 32895
rect 22738 32892 22744 32904
rect 22419 32864 22744 32892
rect 22419 32861 22431 32864
rect 22373 32855 22431 32861
rect 22738 32852 22744 32864
rect 22796 32852 22802 32904
rect 23584 32836 23612 32932
rect 24949 32895 25007 32901
rect 24949 32861 24961 32895
rect 24995 32892 25007 32895
rect 25038 32892 25044 32904
rect 24995 32864 25044 32892
rect 24995 32861 25007 32864
rect 24949 32855 25007 32861
rect 25038 32852 25044 32864
rect 25096 32852 25102 32904
rect 27614 32892 27620 32904
rect 27575 32864 27620 32892
rect 27614 32852 27620 32864
rect 27672 32852 27678 32904
rect 30650 32852 30656 32904
rect 30708 32892 30714 32904
rect 30745 32895 30803 32901
rect 30745 32892 30757 32895
rect 30708 32864 30757 32892
rect 30708 32852 30714 32864
rect 30745 32861 30757 32864
rect 30791 32861 30803 32895
rect 30745 32855 30803 32861
rect 18340 32796 20208 32824
rect 20257 32827 20315 32833
rect 11992 32728 12480 32756
rect 14826 32716 14832 32768
rect 14884 32756 14890 32768
rect 15473 32759 15531 32765
rect 15473 32756 15485 32759
rect 14884 32728 15485 32756
rect 14884 32716 14890 32728
rect 15473 32725 15485 32728
rect 15519 32725 15531 32759
rect 15473 32719 15531 32725
rect 17678 32716 17684 32768
rect 17736 32756 17742 32768
rect 18340 32756 18368 32796
rect 20257 32793 20269 32827
rect 20303 32824 20315 32827
rect 23290 32824 23296 32836
rect 20303 32796 20418 32824
rect 20303 32793 20315 32796
rect 20257 32787 20315 32793
rect 20390 32768 20418 32796
rect 20346 32756 20352 32768
rect 17736 32728 18368 32756
rect 20285 32728 20352 32756
rect 17736 32716 17742 32728
rect 20346 32716 20352 32728
rect 20404 32756 20418 32768
rect 20548 32796 23296 32824
rect 20548 32756 20576 32796
rect 23290 32784 23296 32796
rect 23348 32824 23354 32836
rect 23385 32827 23443 32833
rect 23385 32824 23397 32827
rect 23348 32796 23397 32824
rect 23348 32784 23354 32796
rect 23385 32793 23397 32796
rect 23431 32793 23443 32827
rect 23566 32824 23572 32836
rect 23527 32796 23572 32824
rect 23385 32787 23443 32793
rect 23566 32784 23572 32796
rect 23624 32784 23630 32836
rect 25216 32827 25274 32833
rect 25216 32793 25228 32827
rect 25262 32824 25274 32827
rect 25314 32824 25320 32836
rect 25262 32796 25320 32824
rect 25262 32793 25274 32796
rect 25216 32787 25274 32793
rect 25314 32784 25320 32796
rect 25372 32784 25378 32836
rect 27884 32827 27942 32833
rect 27884 32793 27896 32827
rect 27930 32824 27942 32827
rect 28166 32824 28172 32836
rect 27930 32796 28172 32824
rect 27930 32793 27942 32796
rect 27884 32787 27942 32793
rect 28166 32784 28172 32796
rect 28224 32784 28230 32836
rect 20404 32728 20576 32756
rect 22281 32759 22339 32765
rect 20404 32716 20410 32728
rect 22281 32725 22293 32759
rect 22327 32756 22339 32759
rect 23474 32756 23480 32768
rect 22327 32728 23480 32756
rect 22327 32725 22339 32728
rect 22281 32719 22339 32725
rect 23474 32716 23480 32728
rect 23532 32716 23538 32768
rect 26142 32716 26148 32768
rect 26200 32756 26206 32768
rect 26329 32759 26387 32765
rect 26329 32756 26341 32759
rect 26200 32728 26341 32756
rect 26200 32716 26206 32728
rect 26329 32725 26341 32728
rect 26375 32725 26387 32759
rect 30558 32756 30564 32768
rect 30519 32728 30564 32756
rect 26329 32719 26387 32725
rect 30558 32716 30564 32728
rect 30616 32716 30622 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 10965 32555 11023 32561
rect 10965 32521 10977 32555
rect 11011 32552 11023 32555
rect 11054 32552 11060 32564
rect 11011 32524 11060 32552
rect 11011 32521 11023 32524
rect 10965 32515 11023 32521
rect 11054 32512 11060 32524
rect 11112 32512 11118 32564
rect 15378 32512 15384 32564
rect 15436 32552 15442 32564
rect 16025 32555 16083 32561
rect 16025 32552 16037 32555
rect 15436 32524 16037 32552
rect 15436 32512 15442 32524
rect 16025 32521 16037 32524
rect 16071 32521 16083 32555
rect 20438 32552 20444 32564
rect 16025 32515 16083 32521
rect 16960 32524 19564 32552
rect 20399 32524 20444 32552
rect 9674 32444 9680 32496
rect 9732 32484 9738 32496
rect 9830 32487 9888 32493
rect 9830 32484 9842 32487
rect 9732 32456 9842 32484
rect 9732 32444 9738 32456
rect 9830 32453 9842 32456
rect 9876 32453 9888 32487
rect 9830 32447 9888 32453
rect 10778 32444 10784 32496
rect 10836 32484 10842 32496
rect 11517 32487 11575 32493
rect 11517 32484 11529 32487
rect 10836 32456 11529 32484
rect 10836 32444 10842 32456
rect 11517 32453 11529 32456
rect 11563 32453 11575 32487
rect 11517 32447 11575 32453
rect 12406 32456 14228 32484
rect 5813 32419 5871 32425
rect 5813 32385 5825 32419
rect 5859 32385 5871 32419
rect 5813 32379 5871 32385
rect 5828 32348 5856 32379
rect 5902 32376 5908 32428
rect 5960 32416 5966 32428
rect 6549 32419 6607 32425
rect 6549 32416 6561 32419
rect 5960 32388 6561 32416
rect 5960 32376 5966 32388
rect 6549 32385 6561 32388
rect 6595 32385 6607 32419
rect 6549 32379 6607 32385
rect 7929 32419 7987 32425
rect 7929 32385 7941 32419
rect 7975 32416 7987 32419
rect 8110 32416 8116 32428
rect 7975 32388 8116 32416
rect 7975 32385 7987 32388
rect 7929 32379 7987 32385
rect 8110 32376 8116 32388
rect 8168 32376 8174 32428
rect 11698 32416 11704 32428
rect 11659 32388 11704 32416
rect 11698 32376 11704 32388
rect 11756 32416 11762 32428
rect 12406 32416 12434 32456
rect 11756 32388 12434 32416
rect 11756 32376 11762 32388
rect 13262 32376 13268 32428
rect 13320 32416 13326 32428
rect 13449 32419 13507 32425
rect 13449 32416 13461 32419
rect 13320 32388 13461 32416
rect 13320 32376 13326 32388
rect 13449 32385 13461 32388
rect 13495 32385 13507 32419
rect 13449 32379 13507 32385
rect 6730 32348 6736 32360
rect 5828 32320 6736 32348
rect 6730 32308 6736 32320
rect 6788 32308 6794 32360
rect 9306 32308 9312 32360
rect 9364 32348 9370 32360
rect 9585 32351 9643 32357
rect 9585 32348 9597 32351
rect 9364 32320 9597 32348
rect 9364 32308 9370 32320
rect 9585 32317 9597 32320
rect 9631 32317 9643 32351
rect 9585 32311 9643 32317
rect 11974 32308 11980 32360
rect 12032 32348 12038 32360
rect 12989 32351 13047 32357
rect 12989 32348 13001 32351
rect 12032 32320 13001 32348
rect 12032 32308 12038 32320
rect 12989 32317 13001 32320
rect 13035 32317 13047 32351
rect 12989 32311 13047 32317
rect 13357 32351 13415 32357
rect 13357 32317 13369 32351
rect 13403 32348 13415 32351
rect 13814 32348 13820 32360
rect 13403 32320 13820 32348
rect 13403 32317 13415 32320
rect 13357 32311 13415 32317
rect 13814 32308 13820 32320
rect 13872 32308 13878 32360
rect 14200 32348 14228 32456
rect 14458 32444 14464 32496
rect 14516 32484 14522 32496
rect 14921 32487 14979 32493
rect 14921 32484 14933 32487
rect 14516 32456 14933 32484
rect 14516 32444 14522 32456
rect 14921 32453 14933 32456
rect 14967 32453 14979 32487
rect 14921 32447 14979 32453
rect 15013 32487 15071 32493
rect 15013 32453 15025 32487
rect 15059 32484 15071 32487
rect 15654 32484 15660 32496
rect 15059 32456 15660 32484
rect 15059 32453 15071 32456
rect 15013 32447 15071 32453
rect 15654 32444 15660 32456
rect 15712 32444 15718 32496
rect 14642 32416 14648 32428
rect 14603 32388 14648 32416
rect 14642 32376 14648 32388
rect 14700 32376 14706 32428
rect 14826 32425 14832 32428
rect 14793 32419 14832 32425
rect 14793 32385 14805 32419
rect 14793 32379 14832 32385
rect 14826 32376 14832 32379
rect 14884 32376 14890 32428
rect 15102 32416 15108 32428
rect 15160 32425 15166 32428
rect 15068 32388 15108 32416
rect 15102 32376 15108 32388
rect 15160 32379 15168 32425
rect 15933 32419 15991 32425
rect 15933 32385 15945 32419
rect 15979 32385 15991 32419
rect 16758 32416 16764 32428
rect 16719 32388 16764 32416
rect 15933 32379 15991 32385
rect 15160 32376 15166 32379
rect 15010 32348 15016 32360
rect 14200 32320 15016 32348
rect 15010 32308 15016 32320
rect 15068 32308 15074 32360
rect 15948 32348 15976 32379
rect 16758 32376 16764 32388
rect 16816 32376 16822 32428
rect 16960 32425 16988 32524
rect 17037 32487 17095 32493
rect 17037 32453 17049 32487
rect 17083 32484 17095 32487
rect 17862 32484 17868 32496
rect 17083 32456 17868 32484
rect 17083 32453 17095 32456
rect 17037 32447 17095 32453
rect 17862 32444 17868 32456
rect 17920 32444 17926 32496
rect 18684 32487 18742 32493
rect 18684 32453 18696 32487
rect 18730 32484 18742 32487
rect 19242 32484 19248 32496
rect 18730 32456 19248 32484
rect 18730 32453 18742 32456
rect 18684 32447 18742 32453
rect 19242 32444 19248 32456
rect 19300 32444 19306 32496
rect 19536 32484 19564 32524
rect 20438 32512 20444 32524
rect 20496 32512 20502 32564
rect 22094 32512 22100 32564
rect 22152 32552 22158 32564
rect 22465 32555 22523 32561
rect 22465 32552 22477 32555
rect 22152 32524 22477 32552
rect 22152 32512 22158 32524
rect 22465 32521 22477 32524
rect 22511 32521 22523 32555
rect 22465 32515 22523 32521
rect 22738 32512 22744 32564
rect 22796 32552 22802 32564
rect 23290 32552 23296 32564
rect 22796 32524 23296 32552
rect 22796 32512 22802 32524
rect 23290 32512 23296 32524
rect 23348 32512 23354 32564
rect 23658 32512 23664 32564
rect 23716 32552 23722 32564
rect 24489 32555 24547 32561
rect 24489 32552 24501 32555
rect 23716 32524 24501 32552
rect 23716 32512 23722 32524
rect 24489 32521 24501 32524
rect 24535 32521 24547 32555
rect 25314 32552 25320 32564
rect 25275 32524 25320 32552
rect 24489 32515 24547 32521
rect 25314 32512 25320 32524
rect 25372 32512 25378 32564
rect 25774 32512 25780 32564
rect 25832 32552 25838 32564
rect 27706 32552 27712 32564
rect 25832 32524 27712 32552
rect 25832 32512 25838 32524
rect 27706 32512 27712 32524
rect 27764 32512 27770 32564
rect 28166 32552 28172 32564
rect 28127 32524 28172 32552
rect 28166 32512 28172 32524
rect 28224 32512 28230 32564
rect 28537 32555 28595 32561
rect 28537 32521 28549 32555
rect 28583 32552 28595 32555
rect 28718 32552 28724 32564
rect 28583 32524 28724 32552
rect 28583 32521 28595 32524
rect 28537 32515 28595 32521
rect 28718 32512 28724 32524
rect 28776 32512 28782 32564
rect 31573 32555 31631 32561
rect 31573 32552 31585 32555
rect 28828 32524 31585 32552
rect 28828 32484 28856 32524
rect 31573 32521 31585 32524
rect 31619 32521 31631 32555
rect 31573 32515 31631 32521
rect 19536 32456 28856 32484
rect 30460 32487 30518 32493
rect 30460 32453 30472 32487
rect 30506 32484 30518 32487
rect 30558 32484 30564 32496
rect 30506 32456 30564 32484
rect 30506 32453 30518 32456
rect 30460 32447 30518 32453
rect 30558 32444 30564 32456
rect 30616 32444 30622 32496
rect 16909 32419 16988 32425
rect 16909 32385 16921 32419
rect 16955 32388 16988 32419
rect 16955 32385 16967 32388
rect 16909 32379 16967 32385
rect 17126 32376 17132 32428
rect 17184 32416 17190 32428
rect 17310 32425 17316 32428
rect 17267 32419 17316 32425
rect 17184 32388 17229 32416
rect 17184 32376 17190 32388
rect 17267 32385 17279 32419
rect 17313 32385 17316 32419
rect 17267 32379 17316 32385
rect 17310 32376 17316 32379
rect 17368 32376 17374 32428
rect 20346 32416 20352 32428
rect 20307 32388 20352 32416
rect 20346 32376 20352 32388
rect 20404 32376 20410 32428
rect 24118 32376 24124 32428
rect 24176 32416 24182 32428
rect 24394 32416 24400 32428
rect 24176 32388 24400 32416
rect 24176 32376 24182 32388
rect 24394 32376 24400 32388
rect 24452 32376 24458 32428
rect 24578 32416 24584 32428
rect 24539 32388 24584 32416
rect 24578 32376 24584 32388
rect 24636 32376 24642 32428
rect 25501 32419 25559 32425
rect 25501 32385 25513 32419
rect 25547 32416 25559 32419
rect 25590 32416 25596 32428
rect 25547 32388 25596 32416
rect 25547 32385 25559 32388
rect 25501 32379 25559 32385
rect 25590 32376 25596 32388
rect 25648 32376 25654 32428
rect 25685 32419 25743 32425
rect 25685 32385 25697 32419
rect 25731 32385 25743 32419
rect 25685 32379 25743 32385
rect 16666 32348 16672 32360
rect 15948 32320 16672 32348
rect 16666 32308 16672 32320
rect 16724 32348 16730 32360
rect 17862 32348 17868 32360
rect 16724 32320 17868 32348
rect 16724 32308 16730 32320
rect 17862 32308 17868 32320
rect 17920 32308 17926 32360
rect 18417 32351 18475 32357
rect 18417 32348 18429 32351
rect 17972 32320 18429 32348
rect 15194 32280 15200 32292
rect 10520 32252 15200 32280
rect 5258 32172 5264 32224
rect 5316 32212 5322 32224
rect 5629 32215 5687 32221
rect 5629 32212 5641 32215
rect 5316 32184 5641 32212
rect 5316 32172 5322 32184
rect 5629 32181 5641 32184
rect 5675 32181 5687 32215
rect 6362 32212 6368 32224
rect 6323 32184 6368 32212
rect 5629 32175 5687 32181
rect 6362 32172 6368 32184
rect 6420 32172 6426 32224
rect 7742 32212 7748 32224
rect 7703 32184 7748 32212
rect 7742 32172 7748 32184
rect 7800 32172 7806 32224
rect 9490 32172 9496 32224
rect 9548 32212 9554 32224
rect 10520 32212 10548 32252
rect 15194 32240 15200 32252
rect 15252 32280 15258 32292
rect 15562 32280 15568 32292
rect 15252 32252 15568 32280
rect 15252 32240 15258 32252
rect 15562 32240 15568 32252
rect 15620 32240 15626 32292
rect 9548 32184 10548 32212
rect 9548 32172 9554 32184
rect 11054 32172 11060 32224
rect 11112 32212 11118 32224
rect 11885 32215 11943 32221
rect 11885 32212 11897 32215
rect 11112 32184 11897 32212
rect 11112 32172 11118 32184
rect 11885 32181 11897 32184
rect 11931 32181 11943 32215
rect 13630 32212 13636 32224
rect 13591 32184 13636 32212
rect 11885 32175 11943 32181
rect 13630 32172 13636 32184
rect 13688 32172 13694 32224
rect 15289 32215 15347 32221
rect 15289 32181 15301 32215
rect 15335 32212 15347 32215
rect 15378 32212 15384 32224
rect 15335 32184 15384 32212
rect 15335 32181 15347 32184
rect 15289 32175 15347 32181
rect 15378 32172 15384 32184
rect 15436 32172 15442 32224
rect 16666 32172 16672 32224
rect 16724 32212 16730 32224
rect 17405 32215 17463 32221
rect 17405 32212 17417 32215
rect 16724 32184 17417 32212
rect 16724 32172 16730 32184
rect 17405 32181 17417 32184
rect 17451 32181 17463 32215
rect 17405 32175 17463 32181
rect 17494 32172 17500 32224
rect 17552 32212 17558 32224
rect 17972 32212 18000 32320
rect 18417 32317 18429 32320
rect 18463 32317 18475 32351
rect 18417 32311 18475 32317
rect 20530 32308 20536 32360
rect 20588 32348 20594 32360
rect 21821 32351 21879 32357
rect 21821 32348 21833 32351
rect 20588 32320 21833 32348
rect 20588 32308 20594 32320
rect 21821 32317 21833 32320
rect 21867 32317 21879 32351
rect 21821 32311 21879 32317
rect 22094 32308 22100 32360
rect 22152 32348 22158 32360
rect 22189 32351 22247 32357
rect 22189 32348 22201 32351
rect 22152 32320 22201 32348
rect 22152 32308 22158 32320
rect 22189 32317 22201 32320
rect 22235 32317 22247 32351
rect 22189 32311 22247 32317
rect 22281 32351 22339 32357
rect 22281 32317 22293 32351
rect 22327 32317 22339 32351
rect 22281 32311 22339 32317
rect 19518 32240 19524 32292
rect 19576 32280 19582 32292
rect 19797 32283 19855 32289
rect 19797 32280 19809 32283
rect 19576 32252 19809 32280
rect 19576 32240 19582 32252
rect 19797 32249 19809 32252
rect 19843 32249 19855 32283
rect 19797 32243 19855 32249
rect 20438 32240 20444 32292
rect 20496 32280 20502 32292
rect 22296 32280 22324 32311
rect 25314 32308 25320 32360
rect 25372 32348 25378 32360
rect 25700 32348 25728 32379
rect 25774 32376 25780 32428
rect 25832 32416 25838 32428
rect 27430 32416 27436 32428
rect 25832 32388 25877 32416
rect 27391 32388 27436 32416
rect 25832 32376 25838 32388
rect 27430 32376 27436 32388
rect 27488 32376 27494 32428
rect 27617 32419 27675 32425
rect 27617 32416 27629 32419
rect 27540 32388 27629 32416
rect 26142 32348 26148 32360
rect 25372 32320 26148 32348
rect 25372 32308 25378 32320
rect 26142 32308 26148 32320
rect 26200 32308 26206 32360
rect 25866 32280 25872 32292
rect 20496 32252 25872 32280
rect 20496 32240 20502 32252
rect 25866 32240 25872 32252
rect 25924 32240 25930 32292
rect 27540 32280 27568 32388
rect 27617 32385 27629 32388
rect 27663 32385 27675 32419
rect 27617 32379 27675 32385
rect 27706 32376 27712 32428
rect 27764 32416 27770 32428
rect 28350 32416 28356 32428
rect 27764 32388 27809 32416
rect 28311 32388 28356 32416
rect 27764 32376 27770 32388
rect 28350 32376 28356 32388
rect 28408 32376 28414 32428
rect 28629 32419 28687 32425
rect 28629 32385 28641 32419
rect 28675 32385 28687 32419
rect 28629 32379 28687 32385
rect 27724 32348 27752 32376
rect 28644 32348 28672 32379
rect 30190 32348 30196 32360
rect 27724 32320 28672 32348
rect 30151 32320 30196 32348
rect 30190 32308 30196 32320
rect 30248 32308 30254 32360
rect 28534 32280 28540 32292
rect 27540 32252 28540 32280
rect 28534 32240 28540 32252
rect 28592 32240 28598 32292
rect 17552 32184 18000 32212
rect 17552 32172 17558 32184
rect 18230 32172 18236 32224
rect 18288 32212 18294 32224
rect 24026 32212 24032 32224
rect 18288 32184 24032 32212
rect 18288 32172 18294 32184
rect 24026 32172 24032 32184
rect 24084 32172 24090 32224
rect 27249 32215 27307 32221
rect 27249 32181 27261 32215
rect 27295 32212 27307 32215
rect 27798 32212 27804 32224
rect 27295 32184 27804 32212
rect 27295 32181 27307 32184
rect 27249 32175 27307 32181
rect 27798 32172 27804 32184
rect 27856 32172 27862 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 10597 32011 10655 32017
rect 10597 31977 10609 32011
rect 10643 32008 10655 32011
rect 11698 32008 11704 32020
rect 10643 31980 11704 32008
rect 10643 31977 10655 31980
rect 10597 31971 10655 31977
rect 11698 31968 11704 31980
rect 11756 31968 11762 32020
rect 11974 31968 11980 32020
rect 12032 32008 12038 32020
rect 13541 32011 13599 32017
rect 12032 31980 13492 32008
rect 12032 31968 12038 31980
rect 13464 31940 13492 31980
rect 13541 31977 13553 32011
rect 13587 32008 13599 32011
rect 13814 32008 13820 32020
rect 13587 31980 13820 32008
rect 13587 31977 13599 31980
rect 13541 31971 13599 31977
rect 13814 31968 13820 31980
rect 13872 31968 13878 32020
rect 14182 31968 14188 32020
rect 14240 32008 14246 32020
rect 15194 32008 15200 32020
rect 14240 31980 15200 32008
rect 14240 31968 14246 31980
rect 15194 31968 15200 31980
rect 15252 32008 15258 32020
rect 16945 32011 17003 32017
rect 16945 32008 16957 32011
rect 15252 31980 16957 32008
rect 15252 31968 15258 31980
rect 16945 31977 16957 31980
rect 16991 32008 17003 32011
rect 17310 32008 17316 32020
rect 16991 31980 17316 32008
rect 16991 31977 17003 31980
rect 16945 31971 17003 31977
rect 17310 31968 17316 31980
rect 17368 32008 17374 32020
rect 17494 32008 17500 32020
rect 17368 31980 17500 32008
rect 17368 31968 17374 31980
rect 17494 31968 17500 31980
rect 17552 31968 17558 32020
rect 17972 31980 18920 32008
rect 13464 31912 16712 31940
rect 13630 31832 13636 31884
rect 13688 31872 13694 31884
rect 14734 31872 14740 31884
rect 13688 31844 14320 31872
rect 13688 31832 13694 31844
rect 4982 31804 4988 31816
rect 4895 31776 4988 31804
rect 4982 31764 4988 31776
rect 5040 31804 5046 31816
rect 7006 31804 7012 31816
rect 5040 31776 5396 31804
rect 5040 31764 5046 31776
rect 5258 31745 5264 31748
rect 5252 31736 5264 31745
rect 5219 31708 5264 31736
rect 5252 31699 5264 31708
rect 5258 31696 5264 31699
rect 5316 31696 5322 31748
rect 5368 31736 5396 31776
rect 6886 31776 7012 31804
rect 6886 31748 6914 31776
rect 7006 31764 7012 31776
rect 7064 31764 7070 31816
rect 7276 31807 7334 31813
rect 7276 31773 7288 31807
rect 7322 31804 7334 31807
rect 7742 31804 7748 31816
rect 7322 31776 7748 31804
rect 7322 31773 7334 31776
rect 7276 31767 7334 31773
rect 7742 31764 7748 31776
rect 7800 31764 7806 31816
rect 9030 31764 9036 31816
rect 9088 31804 9094 31816
rect 9217 31807 9275 31813
rect 9217 31804 9229 31807
rect 9088 31776 9229 31804
rect 9088 31764 9094 31776
rect 9217 31773 9229 31776
rect 9263 31804 9275 31807
rect 9306 31804 9312 31816
rect 9263 31776 9312 31804
rect 9263 31773 9275 31776
rect 9217 31767 9275 31773
rect 9306 31764 9312 31776
rect 9364 31804 9370 31816
rect 14292 31813 14320 31844
rect 14476 31844 14740 31872
rect 14476 31813 14504 31844
rect 14734 31832 14740 31844
rect 14792 31832 14798 31884
rect 16684 31872 16712 31912
rect 16758 31900 16764 31952
rect 16816 31940 16822 31952
rect 17865 31943 17923 31949
rect 17865 31940 17877 31943
rect 16816 31912 17877 31940
rect 16816 31900 16822 31912
rect 17865 31909 17877 31912
rect 17911 31909 17923 31943
rect 17865 31903 17923 31909
rect 17972 31872 18000 31980
rect 18230 31940 18236 31952
rect 16684 31844 18000 31872
rect 18156 31912 18236 31940
rect 12161 31807 12219 31813
rect 12161 31804 12173 31807
rect 9364 31776 12173 31804
rect 9364 31764 9370 31776
rect 12161 31773 12173 31776
rect 12207 31773 12219 31807
rect 12161 31767 12219 31773
rect 12428 31807 12486 31813
rect 12428 31773 12440 31807
rect 12474 31804 12486 31807
rect 14093 31807 14151 31813
rect 14093 31804 14105 31807
rect 12474 31776 14105 31804
rect 12474 31773 12486 31776
rect 12428 31767 12486 31773
rect 14093 31773 14105 31776
rect 14139 31773 14151 31807
rect 14093 31767 14151 31773
rect 14277 31807 14335 31813
rect 14277 31773 14289 31807
rect 14323 31773 14335 31807
rect 14277 31767 14335 31773
rect 14461 31807 14519 31813
rect 14461 31773 14473 31807
rect 14507 31773 14519 31807
rect 14461 31767 14519 31773
rect 14553 31807 14611 31813
rect 14553 31773 14565 31807
rect 14599 31804 14611 31807
rect 14642 31804 14648 31816
rect 14599 31776 14648 31804
rect 14599 31773 14611 31776
rect 14553 31767 14611 31773
rect 14642 31764 14648 31776
rect 14700 31764 14706 31816
rect 15562 31764 15568 31816
rect 15620 31804 15626 31816
rect 15657 31807 15715 31813
rect 15657 31804 15669 31807
rect 15620 31776 15669 31804
rect 15620 31764 15626 31776
rect 15657 31773 15669 31776
rect 15703 31773 15715 31807
rect 18046 31804 18052 31816
rect 18007 31776 18052 31804
rect 15657 31767 15715 31773
rect 18046 31764 18052 31776
rect 18104 31764 18110 31816
rect 18156 31813 18184 31912
rect 18230 31900 18236 31912
rect 18288 31900 18294 31952
rect 18782 31872 18788 31884
rect 18248 31844 18788 31872
rect 18248 31813 18276 31844
rect 18782 31832 18788 31844
rect 18840 31832 18846 31884
rect 18892 31872 18920 31980
rect 19426 31968 19432 32020
rect 19484 32008 19490 32020
rect 19889 32011 19947 32017
rect 19889 32008 19901 32011
rect 19484 31980 19901 32008
rect 19484 31968 19490 31980
rect 19889 31977 19901 31980
rect 19935 31977 19947 32011
rect 19889 31971 19947 31977
rect 23566 31968 23572 32020
rect 23624 32008 23630 32020
rect 24026 32008 24032 32020
rect 23624 31980 24032 32008
rect 23624 31968 23630 31980
rect 24026 31968 24032 31980
rect 24084 31968 24090 32020
rect 25590 31968 25596 32020
rect 25648 32008 25654 32020
rect 26053 32011 26111 32017
rect 26053 32008 26065 32011
rect 25648 31980 26065 32008
rect 25648 31968 25654 31980
rect 26053 31977 26065 31980
rect 26099 31977 26111 32011
rect 26053 31971 26111 31977
rect 27430 31968 27436 32020
rect 27488 32008 27494 32020
rect 28077 32011 28135 32017
rect 28077 32008 28089 32011
rect 27488 31980 28089 32008
rect 27488 31968 27494 31980
rect 28077 31977 28089 31980
rect 28123 31977 28135 32011
rect 30466 32008 30472 32020
rect 30427 31980 30472 32008
rect 28077 31971 28135 31977
rect 30466 31968 30472 31980
rect 30524 31968 30530 32020
rect 30650 32008 30656 32020
rect 30611 31980 30656 32008
rect 30650 31968 30656 31980
rect 30708 31968 30714 32020
rect 22002 31940 22008 31952
rect 21963 31912 22008 31940
rect 22002 31900 22008 31912
rect 22060 31900 22066 31952
rect 29638 31900 29644 31952
rect 29696 31940 29702 31952
rect 30101 31943 30159 31949
rect 30101 31940 30113 31943
rect 29696 31912 30113 31940
rect 29696 31900 29702 31912
rect 30101 31909 30113 31912
rect 30147 31940 30159 31943
rect 31113 31943 31171 31949
rect 31113 31940 31125 31943
rect 30147 31912 31125 31940
rect 30147 31909 30159 31912
rect 30101 31903 30159 31909
rect 31113 31909 31125 31912
rect 31159 31909 31171 31943
rect 31113 31903 31171 31909
rect 19245 31875 19303 31881
rect 19245 31872 19257 31875
rect 18892 31844 19257 31872
rect 19245 31841 19257 31844
rect 19291 31872 19303 31875
rect 20530 31872 20536 31884
rect 19291 31844 20536 31872
rect 19291 31841 19303 31844
rect 19245 31835 19303 31841
rect 20530 31832 20536 31844
rect 20588 31832 20594 31884
rect 22186 31872 22192 31884
rect 22066 31844 22192 31872
rect 18141 31807 18199 31813
rect 18141 31773 18153 31807
rect 18187 31773 18199 31807
rect 18141 31767 18199 31773
rect 18233 31807 18291 31813
rect 18233 31773 18245 31807
rect 18279 31773 18291 31807
rect 18351 31807 18409 31813
rect 18351 31804 18363 31807
rect 18233 31767 18291 31773
rect 18340 31773 18363 31804
rect 18397 31773 18409 31807
rect 18340 31767 18409 31773
rect 18509 31807 18567 31813
rect 18509 31773 18521 31807
rect 18555 31804 18567 31807
rect 18690 31804 18696 31816
rect 18555 31776 18696 31804
rect 18555 31773 18567 31776
rect 18509 31767 18567 31773
rect 6822 31736 6828 31748
rect 5368 31708 6828 31736
rect 6822 31696 6828 31708
rect 6880 31708 6914 31748
rect 9484 31739 9542 31745
rect 6880 31696 6886 31708
rect 9484 31705 9496 31739
rect 9530 31736 9542 31739
rect 9582 31736 9588 31748
rect 9530 31708 9588 31736
rect 9530 31705 9542 31708
rect 9484 31699 9542 31705
rect 9582 31696 9588 31708
rect 9640 31696 9646 31748
rect 17770 31696 17776 31748
rect 17828 31736 17834 31748
rect 17954 31736 17960 31748
rect 17828 31708 17960 31736
rect 17828 31696 17834 31708
rect 17954 31696 17960 31708
rect 18012 31696 18018 31748
rect 6362 31668 6368 31680
rect 6323 31640 6368 31668
rect 6362 31628 6368 31640
rect 6420 31628 6426 31680
rect 8386 31668 8392 31680
rect 8347 31640 8392 31668
rect 8386 31628 8392 31640
rect 8444 31628 8450 31680
rect 8938 31628 8944 31680
rect 8996 31668 9002 31680
rect 13630 31668 13636 31680
rect 8996 31640 13636 31668
rect 8996 31628 9002 31640
rect 13630 31628 13636 31640
rect 13688 31628 13694 31680
rect 18138 31628 18144 31680
rect 18196 31668 18202 31680
rect 18340 31668 18368 31767
rect 18690 31764 18696 31776
rect 18748 31764 18754 31816
rect 19334 31764 19340 31816
rect 19392 31804 19398 31816
rect 19613 31807 19671 31813
rect 19613 31804 19625 31807
rect 19392 31776 19625 31804
rect 19392 31764 19398 31776
rect 19613 31773 19625 31776
rect 19659 31773 19671 31807
rect 19613 31767 19671 31773
rect 19705 31807 19763 31813
rect 19705 31773 19717 31807
rect 19751 31804 19763 31807
rect 20438 31804 20444 31816
rect 19751 31776 20444 31804
rect 19751 31773 19763 31776
rect 19705 31767 19763 31773
rect 19426 31696 19432 31748
rect 19484 31736 19490 31748
rect 19720 31736 19748 31767
rect 20438 31764 20444 31776
rect 20496 31764 20502 31816
rect 20625 31807 20683 31813
rect 20625 31773 20637 31807
rect 20671 31804 20683 31807
rect 22066 31804 22094 31844
rect 22186 31832 22192 31844
rect 22244 31872 22250 31884
rect 22465 31875 22523 31881
rect 22465 31872 22477 31875
rect 22244 31844 22477 31872
rect 22244 31832 22250 31844
rect 22465 31841 22477 31844
rect 22511 31841 22523 31875
rect 25866 31872 25872 31884
rect 25827 31844 25872 31872
rect 22465 31835 22523 31841
rect 25866 31832 25872 31844
rect 25924 31832 25930 31884
rect 27798 31872 27804 31884
rect 27759 31844 27804 31872
rect 27798 31832 27804 31844
rect 27856 31832 27862 31884
rect 20671 31776 22094 31804
rect 25777 31807 25835 31813
rect 20671 31773 20683 31776
rect 20625 31767 20683 31773
rect 25777 31773 25789 31807
rect 25823 31773 25835 31807
rect 25884 31804 25912 31832
rect 27893 31807 27951 31813
rect 27893 31804 27905 31807
rect 25884 31776 27905 31804
rect 25777 31767 25835 31773
rect 27893 31773 27905 31776
rect 27939 31804 27951 31807
rect 27982 31804 27988 31816
rect 27939 31776 27988 31804
rect 27939 31773 27951 31776
rect 27893 31767 27951 31773
rect 20898 31745 20904 31748
rect 19484 31708 19748 31736
rect 19484 31696 19490 31708
rect 20892 31699 20904 31745
rect 20956 31736 20962 31748
rect 20956 31708 20992 31736
rect 20898 31696 20904 31699
rect 20956 31696 20962 31708
rect 21174 31696 21180 31748
rect 21232 31736 21238 31748
rect 21726 31736 21732 31748
rect 21232 31708 21732 31736
rect 21232 31696 21238 31708
rect 21726 31696 21732 31708
rect 21784 31736 21790 31748
rect 22094 31736 22100 31748
rect 21784 31708 22100 31736
rect 21784 31696 21790 31708
rect 22094 31696 22100 31708
rect 22152 31696 22158 31748
rect 22732 31739 22790 31745
rect 22732 31705 22744 31739
rect 22778 31736 22790 31739
rect 23106 31736 23112 31748
rect 22778 31708 23112 31736
rect 22778 31705 22790 31708
rect 22732 31699 22790 31705
rect 23106 31696 23112 31708
rect 23164 31696 23170 31748
rect 24118 31696 24124 31748
rect 24176 31736 24182 31748
rect 25792 31736 25820 31767
rect 27982 31764 27988 31776
rect 28040 31764 28046 31816
rect 30742 31764 30748 31816
rect 30800 31804 30806 31816
rect 31113 31807 31171 31813
rect 31113 31804 31125 31807
rect 30800 31776 31125 31804
rect 30800 31764 30806 31776
rect 31113 31773 31125 31776
rect 31159 31773 31171 31807
rect 31294 31804 31300 31816
rect 31255 31776 31300 31804
rect 31113 31767 31171 31773
rect 31294 31764 31300 31776
rect 31352 31764 31358 31816
rect 24176 31708 25820 31736
rect 24176 31696 24182 31708
rect 18196 31640 18368 31668
rect 18196 31628 18202 31640
rect 23658 31628 23664 31680
rect 23716 31668 23722 31680
rect 23845 31671 23903 31677
rect 23845 31668 23857 31671
rect 23716 31640 23857 31668
rect 23716 31628 23722 31640
rect 23845 31637 23857 31640
rect 23891 31668 23903 31671
rect 24394 31668 24400 31680
rect 23891 31640 24400 31668
rect 23891 31637 23903 31640
rect 23845 31631 23903 31637
rect 24394 31628 24400 31640
rect 24452 31628 24458 31680
rect 25406 31668 25412 31680
rect 25367 31640 25412 31668
rect 25406 31628 25412 31640
rect 25464 31668 25470 31680
rect 27433 31671 27491 31677
rect 27433 31668 27445 31671
rect 25464 31640 27445 31668
rect 25464 31628 25470 31640
rect 27433 31637 27445 31640
rect 27479 31668 27491 31671
rect 27522 31668 27528 31680
rect 27479 31640 27528 31668
rect 27479 31637 27491 31640
rect 27433 31631 27491 31637
rect 27522 31628 27528 31640
rect 27580 31628 27586 31680
rect 30466 31668 30472 31680
rect 30427 31640 30472 31668
rect 30466 31628 30472 31640
rect 30524 31628 30530 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 5813 31467 5871 31473
rect 5813 31433 5825 31467
rect 5859 31464 5871 31467
rect 5902 31464 5908 31476
rect 5859 31436 5908 31464
rect 5859 31433 5871 31436
rect 5813 31427 5871 31433
rect 5902 31424 5908 31436
rect 5960 31424 5966 31476
rect 6546 31464 6552 31476
rect 6604 31473 6610 31476
rect 6604 31467 6623 31473
rect 6288 31436 6552 31464
rect 5445 31399 5503 31405
rect 5445 31365 5457 31399
rect 5491 31365 5503 31399
rect 5445 31359 5503 31365
rect 5661 31399 5719 31405
rect 5661 31365 5673 31399
rect 5707 31396 5719 31399
rect 6288 31396 6316 31436
rect 6546 31424 6552 31436
rect 6611 31433 6623 31467
rect 6730 31464 6736 31476
rect 6691 31436 6736 31464
rect 6604 31427 6623 31433
rect 6604 31424 6610 31427
rect 6730 31424 6736 31436
rect 6788 31424 6794 31476
rect 9582 31464 9588 31476
rect 9543 31436 9588 31464
rect 9582 31424 9588 31436
rect 9640 31424 9646 31476
rect 9950 31424 9956 31476
rect 10008 31424 10014 31476
rect 12802 31424 12808 31476
rect 12860 31464 12866 31476
rect 12897 31467 12955 31473
rect 12897 31464 12909 31467
rect 12860 31436 12909 31464
rect 12860 31424 12866 31436
rect 12897 31433 12909 31436
rect 12943 31433 12955 31467
rect 12897 31427 12955 31433
rect 13630 31424 13636 31476
rect 13688 31464 13694 31476
rect 13725 31467 13783 31473
rect 13725 31464 13737 31467
rect 13688 31436 13737 31464
rect 13688 31424 13694 31436
rect 13725 31433 13737 31436
rect 13771 31433 13783 31467
rect 13725 31427 13783 31433
rect 13814 31424 13820 31476
rect 13872 31464 13878 31476
rect 14642 31464 14648 31476
rect 13872 31436 14648 31464
rect 13872 31424 13878 31436
rect 14642 31424 14648 31436
rect 14700 31464 14706 31476
rect 18230 31464 18236 31476
rect 14700 31436 18236 31464
rect 14700 31424 14706 31436
rect 18230 31424 18236 31436
rect 18288 31424 18294 31476
rect 20809 31467 20867 31473
rect 20809 31433 20821 31467
rect 20855 31464 20867 31467
rect 20898 31464 20904 31476
rect 20855 31436 20904 31464
rect 20855 31433 20867 31436
rect 20809 31427 20867 31433
rect 20898 31424 20904 31436
rect 20956 31424 20962 31476
rect 21174 31464 21180 31476
rect 21135 31436 21180 31464
rect 21174 31424 21180 31436
rect 21232 31424 21238 31476
rect 21818 31464 21824 31476
rect 21731 31436 21824 31464
rect 21818 31424 21824 31436
rect 21876 31464 21882 31476
rect 27522 31464 27528 31476
rect 21876 31436 23244 31464
rect 27483 31436 27528 31464
rect 21876 31424 21882 31436
rect 5707 31368 6316 31396
rect 6365 31399 6423 31405
rect 5707 31365 5719 31368
rect 5661 31359 5719 31365
rect 6365 31365 6377 31399
rect 6411 31365 6423 31399
rect 6365 31359 6423 31365
rect 5460 31328 5488 31359
rect 6380 31328 6408 31359
rect 6730 31328 6736 31340
rect 5460 31300 6736 31328
rect 6730 31288 6736 31300
rect 6788 31288 6794 31340
rect 7006 31288 7012 31340
rect 7064 31328 7070 31340
rect 7193 31331 7251 31337
rect 7193 31328 7205 31331
rect 7064 31300 7205 31328
rect 7064 31288 7070 31300
rect 7193 31297 7205 31300
rect 7239 31297 7251 31331
rect 7193 31291 7251 31297
rect 7282 31288 7288 31340
rect 7340 31328 7346 31340
rect 7449 31331 7507 31337
rect 7449 31328 7461 31331
rect 7340 31300 7461 31328
rect 7340 31288 7346 31300
rect 7449 31297 7461 31300
rect 7495 31297 7507 31331
rect 7449 31291 7507 31297
rect 9674 31288 9680 31340
rect 9732 31328 9738 31340
rect 9968 31337 9996 31424
rect 11532 31368 14228 31396
rect 9861 31331 9919 31337
rect 9861 31328 9873 31331
rect 9732 31300 9873 31328
rect 9732 31288 9738 31300
rect 9861 31297 9873 31300
rect 9907 31297 9919 31331
rect 9861 31291 9919 31297
rect 9953 31331 10011 31337
rect 9953 31297 9965 31331
rect 9999 31297 10011 31331
rect 9953 31291 10011 31297
rect 10045 31331 10103 31337
rect 10045 31297 10057 31331
rect 10091 31297 10103 31331
rect 10226 31328 10232 31340
rect 10187 31300 10232 31328
rect 10045 31291 10103 31297
rect 10060 31260 10088 31291
rect 10226 31288 10232 31300
rect 10284 31288 10290 31340
rect 11532 31337 11560 31368
rect 14200 31340 14228 31368
rect 16482 31356 16488 31408
rect 16540 31396 16546 31408
rect 16669 31399 16727 31405
rect 16669 31396 16681 31399
rect 16540 31368 16681 31396
rect 16540 31356 16546 31368
rect 16669 31365 16681 31368
rect 16715 31396 16727 31399
rect 18506 31396 18512 31408
rect 16715 31368 18512 31396
rect 16715 31365 16727 31368
rect 16669 31359 16727 31365
rect 18506 31356 18512 31368
rect 18564 31396 18570 31408
rect 18690 31396 18696 31408
rect 18564 31368 18696 31396
rect 18564 31356 18570 31368
rect 18690 31356 18696 31368
rect 18748 31396 18754 31408
rect 19061 31399 19119 31405
rect 19061 31396 19073 31399
rect 18748 31368 19073 31396
rect 18748 31356 18754 31368
rect 19061 31365 19073 31368
rect 19107 31365 19119 31399
rect 19061 31359 19119 31365
rect 19245 31399 19303 31405
rect 19245 31365 19257 31399
rect 19291 31396 19303 31399
rect 19426 31396 19432 31408
rect 19291 31368 19432 31396
rect 19291 31365 19303 31368
rect 19245 31359 19303 31365
rect 19426 31356 19432 31368
rect 19484 31356 19490 31408
rect 23216 31405 23244 31436
rect 27522 31424 27528 31436
rect 27580 31424 27586 31476
rect 28169 31467 28227 31473
rect 28169 31433 28181 31467
rect 28215 31464 28227 31467
rect 28350 31464 28356 31476
rect 28215 31436 28356 31464
rect 28215 31433 28227 31436
rect 28169 31427 28227 31433
rect 28350 31424 28356 31436
rect 28408 31424 28414 31476
rect 30466 31424 30472 31476
rect 30524 31464 30530 31476
rect 30837 31467 30895 31473
rect 30837 31464 30849 31467
rect 30524 31436 30849 31464
rect 30524 31424 30530 31436
rect 30837 31433 30849 31436
rect 30883 31433 30895 31467
rect 30837 31427 30895 31433
rect 22465 31399 22523 31405
rect 22465 31396 22477 31399
rect 21008 31368 22477 31396
rect 11517 31331 11575 31337
rect 11517 31297 11529 31331
rect 11563 31297 11575 31331
rect 11517 31291 11575 31297
rect 11784 31331 11842 31337
rect 11784 31297 11796 31331
rect 11830 31328 11842 31331
rect 13357 31331 13415 31337
rect 13357 31328 13369 31331
rect 11830 31300 13369 31328
rect 11830 31297 11842 31300
rect 11784 31291 11842 31297
rect 13357 31297 13369 31300
rect 13403 31297 13415 31331
rect 13538 31328 13544 31340
rect 13499 31300 13544 31328
rect 13357 31291 13415 31297
rect 13538 31288 13544 31300
rect 13596 31288 13602 31340
rect 13814 31328 13820 31340
rect 13775 31300 13820 31328
rect 13814 31288 13820 31300
rect 13872 31288 13878 31340
rect 14182 31288 14188 31340
rect 14240 31328 14246 31340
rect 14277 31331 14335 31337
rect 14277 31328 14289 31331
rect 14240 31300 14289 31328
rect 14240 31288 14246 31300
rect 14277 31297 14289 31300
rect 14323 31297 14335 31331
rect 14277 31291 14335 31297
rect 14366 31288 14372 31340
rect 14424 31328 14430 31340
rect 14533 31331 14591 31337
rect 14533 31328 14545 31331
rect 14424 31300 14545 31328
rect 14424 31288 14430 31300
rect 14533 31297 14545 31300
rect 14579 31297 14591 31331
rect 16850 31328 16856 31340
rect 16811 31300 16856 31328
rect 14533 31291 14591 31297
rect 16850 31288 16856 31300
rect 16908 31328 16914 31340
rect 17126 31328 17132 31340
rect 16908 31300 17132 31328
rect 16908 31288 16914 31300
rect 17126 31288 17132 31300
rect 17184 31288 17190 31340
rect 18138 31328 18144 31340
rect 18099 31300 18144 31328
rect 18138 31288 18144 31300
rect 18196 31288 18202 31340
rect 20165 31331 20223 31337
rect 20165 31297 20177 31331
rect 20211 31328 20223 31331
rect 20806 31328 20812 31340
rect 20211 31300 20812 31328
rect 20211 31297 20223 31300
rect 20165 31291 20223 31297
rect 20806 31288 20812 31300
rect 20864 31288 20870 31340
rect 21008 31337 21036 31368
rect 22465 31365 22477 31368
rect 22511 31365 22523 31399
rect 22465 31359 22523 31365
rect 23201 31399 23259 31405
rect 23201 31365 23213 31399
rect 23247 31396 23259 31399
rect 24210 31396 24216 31408
rect 23247 31368 24216 31396
rect 23247 31365 23259 31368
rect 23201 31359 23259 31365
rect 24210 31356 24216 31368
rect 24268 31356 24274 31408
rect 28994 31396 29000 31408
rect 24872 31368 29000 31396
rect 20993 31331 21051 31337
rect 20993 31297 21005 31331
rect 21039 31297 21051 31331
rect 20993 31291 21051 31297
rect 21269 31331 21327 31337
rect 21269 31297 21281 31331
rect 21315 31328 21327 31331
rect 22094 31328 22100 31340
rect 21315 31300 22100 31328
rect 21315 31297 21327 31300
rect 21269 31291 21327 31297
rect 11054 31260 11060 31272
rect 10060 31232 11060 31260
rect 11054 31220 11060 31232
rect 11112 31220 11118 31272
rect 18230 31220 18236 31272
rect 18288 31260 18294 31272
rect 21284 31260 21312 31291
rect 22094 31288 22100 31300
rect 22152 31288 22158 31340
rect 22278 31328 22284 31340
rect 22191 31300 22284 31328
rect 22278 31288 22284 31300
rect 22336 31328 22342 31340
rect 23661 31331 23719 31337
rect 23661 31328 23673 31331
rect 22336 31300 23673 31328
rect 22336 31288 22342 31300
rect 23661 31297 23673 31300
rect 23707 31297 23719 31331
rect 23661 31291 23719 31297
rect 18288 31232 21312 31260
rect 18288 31220 18294 31232
rect 22002 31220 22008 31272
rect 22060 31260 22066 31272
rect 22189 31263 22247 31269
rect 22189 31260 22201 31263
rect 22060 31232 22201 31260
rect 22060 31220 22066 31232
rect 22189 31229 22201 31232
rect 22235 31229 22247 31263
rect 23566 31260 23572 31272
rect 23527 31232 23572 31260
rect 22189 31223 22247 31229
rect 23566 31220 23572 31232
rect 23624 31220 23630 31272
rect 18322 31192 18328 31204
rect 18235 31164 18328 31192
rect 18322 31152 18328 31164
rect 18380 31192 18386 31204
rect 24872 31192 24900 31368
rect 28994 31356 29000 31368
rect 29052 31356 29058 31408
rect 30098 31396 30104 31408
rect 29104 31368 30104 31396
rect 24949 31331 25007 31337
rect 24949 31297 24961 31331
rect 24995 31328 25007 31331
rect 25038 31328 25044 31340
rect 24995 31300 25044 31328
rect 24995 31297 25007 31300
rect 24949 31291 25007 31297
rect 25038 31288 25044 31300
rect 25096 31288 25102 31340
rect 25222 31337 25228 31340
rect 25216 31291 25228 31337
rect 25280 31328 25286 31340
rect 27982 31328 27988 31340
rect 25280 31300 25316 31328
rect 27943 31300 27988 31328
rect 25222 31288 25228 31291
rect 25280 31288 25286 31300
rect 27982 31288 27988 31300
rect 28040 31288 28046 31340
rect 28905 31331 28963 31337
rect 28905 31297 28917 31331
rect 28951 31328 28963 31331
rect 29104 31328 29132 31368
rect 30098 31356 30104 31368
rect 30156 31356 30162 31408
rect 29178 31337 29184 31340
rect 28951 31300 29132 31328
rect 28951 31297 28963 31300
rect 28905 31291 28963 31297
rect 29172 31291 29184 31337
rect 29236 31328 29242 31340
rect 30742 31328 30748 31340
rect 29236 31300 29272 31328
rect 30300 31300 30748 31328
rect 29178 31288 29184 31291
rect 29236 31288 29242 31300
rect 27893 31263 27951 31269
rect 27893 31229 27905 31263
rect 27939 31229 27951 31263
rect 27893 31223 27951 31229
rect 18380 31164 24900 31192
rect 27908 31192 27936 31223
rect 27982 31192 27988 31204
rect 27908 31164 27988 31192
rect 18380 31152 18386 31164
rect 27982 31152 27988 31164
rect 28040 31152 28046 31204
rect 5626 31124 5632 31136
rect 5587 31096 5632 31124
rect 5626 31084 5632 31096
rect 5684 31084 5690 31136
rect 6362 31084 6368 31136
rect 6420 31124 6426 31136
rect 6549 31127 6607 31133
rect 6549 31124 6561 31127
rect 6420 31096 6561 31124
rect 6420 31084 6426 31096
rect 6549 31093 6561 31096
rect 6595 31093 6607 31127
rect 8570 31124 8576 31136
rect 8531 31096 8576 31124
rect 6549 31087 6607 31093
rect 8570 31084 8576 31096
rect 8628 31084 8634 31136
rect 15654 31124 15660 31136
rect 15615 31096 15660 31124
rect 15654 31084 15660 31096
rect 15712 31084 15718 31136
rect 17037 31127 17095 31133
rect 17037 31093 17049 31127
rect 17083 31124 17095 31127
rect 17126 31124 17132 31136
rect 17083 31096 17132 31124
rect 17083 31093 17095 31096
rect 17037 31087 17095 31093
rect 17126 31084 17132 31096
rect 17184 31084 17190 31136
rect 17218 31084 17224 31136
rect 17276 31124 17282 31136
rect 20257 31127 20315 31133
rect 20257 31124 20269 31127
rect 17276 31096 20269 31124
rect 17276 31084 17282 31096
rect 20257 31093 20269 31096
rect 20303 31124 20315 31127
rect 20346 31124 20352 31136
rect 20303 31096 20352 31124
rect 20303 31093 20315 31096
rect 20257 31087 20315 31093
rect 20346 31084 20352 31096
rect 20404 31084 20410 31136
rect 23290 31084 23296 31136
rect 23348 31124 23354 31136
rect 23845 31127 23903 31133
rect 23845 31124 23857 31127
rect 23348 31096 23857 31124
rect 23348 31084 23354 31096
rect 23845 31093 23857 31096
rect 23891 31093 23903 31127
rect 23845 31087 23903 31093
rect 26142 31084 26148 31136
rect 26200 31124 26206 31136
rect 26329 31127 26387 31133
rect 26329 31124 26341 31127
rect 26200 31096 26341 31124
rect 26200 31084 26206 31096
rect 26329 31093 26341 31096
rect 26375 31093 26387 31127
rect 26329 31087 26387 31093
rect 28626 31084 28632 31136
rect 28684 31124 28690 31136
rect 30300 31133 30328 31300
rect 30742 31288 30748 31300
rect 30800 31288 30806 31340
rect 30929 31331 30987 31337
rect 30929 31297 30941 31331
rect 30975 31328 30987 31331
rect 31294 31328 31300 31340
rect 30975 31300 31300 31328
rect 30975 31297 30987 31300
rect 30929 31291 30987 31297
rect 31294 31288 31300 31300
rect 31352 31288 31358 31340
rect 30285 31127 30343 31133
rect 30285 31124 30297 31127
rect 28684 31096 30297 31124
rect 28684 31084 28690 31096
rect 30285 31093 30297 31096
rect 30331 31093 30343 31127
rect 30285 31087 30343 31093
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 5626 30880 5632 30932
rect 5684 30920 5690 30932
rect 6365 30923 6423 30929
rect 6365 30920 6377 30923
rect 5684 30892 6377 30920
rect 5684 30880 5690 30892
rect 6365 30889 6377 30892
rect 6411 30889 6423 30923
rect 6365 30883 6423 30889
rect 7101 30923 7159 30929
rect 7101 30889 7113 30923
rect 7147 30920 7159 30923
rect 7282 30920 7288 30932
rect 7147 30892 7288 30920
rect 7147 30889 7159 30892
rect 7101 30883 7159 30889
rect 7282 30880 7288 30892
rect 7340 30880 7346 30932
rect 7929 30923 7987 30929
rect 7929 30889 7941 30923
rect 7975 30889 7987 30923
rect 8110 30920 8116 30932
rect 8071 30892 8116 30920
rect 7929 30883 7987 30889
rect 7944 30852 7972 30883
rect 8110 30880 8116 30892
rect 8168 30880 8174 30932
rect 12713 30923 12771 30929
rect 12713 30889 12725 30923
rect 12759 30920 12771 30923
rect 13538 30920 13544 30932
rect 12759 30892 13544 30920
rect 12759 30889 12771 30892
rect 12713 30883 12771 30889
rect 13538 30880 13544 30892
rect 13596 30880 13602 30932
rect 13630 30880 13636 30932
rect 13688 30880 13694 30932
rect 14093 30923 14151 30929
rect 14093 30889 14105 30923
rect 14139 30920 14151 30923
rect 14366 30920 14372 30932
rect 14139 30892 14372 30920
rect 14139 30889 14151 30892
rect 14093 30883 14151 30889
rect 14366 30880 14372 30892
rect 14424 30880 14430 30932
rect 16114 30880 16120 30932
rect 16172 30920 16178 30932
rect 18782 30920 18788 30932
rect 16172 30892 18788 30920
rect 16172 30880 16178 30892
rect 18782 30880 18788 30892
rect 18840 30880 18846 30932
rect 23106 30920 23112 30932
rect 23067 30892 23112 30920
rect 23106 30880 23112 30892
rect 23164 30880 23170 30932
rect 24489 30923 24547 30929
rect 24489 30889 24501 30923
rect 24535 30920 24547 30923
rect 25222 30920 25228 30932
rect 24535 30892 25228 30920
rect 24535 30889 24547 30892
rect 24489 30883 24547 30889
rect 25222 30880 25228 30892
rect 25280 30880 25286 30932
rect 8386 30852 8392 30864
rect 7944 30824 8392 30852
rect 8386 30812 8392 30824
rect 8444 30812 8450 30864
rect 13648 30852 13676 30880
rect 13556 30824 13676 30852
rect 18693 30855 18751 30861
rect 13556 30796 13584 30824
rect 18693 30821 18705 30855
rect 18739 30852 18751 30855
rect 19150 30852 19156 30864
rect 18739 30824 19156 30852
rect 18739 30821 18751 30824
rect 18693 30815 18751 30821
rect 19150 30812 19156 30824
rect 19208 30852 19214 30864
rect 19208 30824 19334 30852
rect 19208 30812 19214 30824
rect 4982 30784 4988 30796
rect 4943 30756 4988 30784
rect 4982 30744 4988 30756
rect 5040 30744 5046 30796
rect 11974 30744 11980 30796
rect 12032 30784 12038 30796
rect 12069 30787 12127 30793
rect 12069 30784 12081 30787
rect 12032 30756 12081 30784
rect 12032 30744 12038 30756
rect 12069 30753 12081 30756
rect 12115 30753 12127 30787
rect 12069 30747 12127 30753
rect 12437 30787 12495 30793
rect 12437 30753 12449 30787
rect 12483 30784 12495 30787
rect 12802 30784 12808 30796
rect 12483 30756 12808 30784
rect 12483 30753 12495 30756
rect 12437 30747 12495 30753
rect 12802 30744 12808 30756
rect 12860 30744 12866 30796
rect 13538 30744 13544 30796
rect 13596 30744 13602 30796
rect 13630 30744 13636 30796
rect 13688 30784 13694 30796
rect 13688 30756 14872 30784
rect 13688 30744 13694 30756
rect 5252 30719 5310 30725
rect 5252 30685 5264 30719
rect 5298 30716 5310 30719
rect 6270 30716 6276 30728
rect 5298 30688 6276 30716
rect 5298 30685 5310 30688
rect 5252 30679 5310 30685
rect 6270 30676 6276 30688
rect 6328 30676 6334 30728
rect 7282 30716 7288 30728
rect 7243 30688 7288 30716
rect 7282 30676 7288 30688
rect 7340 30676 7346 30728
rect 12529 30719 12587 30725
rect 12529 30685 12541 30719
rect 12575 30716 12587 30719
rect 13262 30716 13268 30728
rect 12575 30688 13268 30716
rect 12575 30685 12587 30688
rect 12529 30679 12587 30685
rect 13262 30676 13268 30688
rect 13320 30716 13326 30728
rect 13648 30716 13676 30744
rect 13320 30688 13676 30716
rect 14369 30719 14427 30725
rect 13320 30676 13326 30688
rect 14369 30685 14381 30719
rect 14415 30685 14427 30719
rect 14369 30679 14427 30685
rect 14461 30719 14519 30725
rect 14461 30685 14473 30719
rect 14507 30685 14519 30719
rect 14461 30679 14519 30685
rect 14553 30719 14611 30725
rect 14553 30685 14565 30719
rect 14599 30685 14611 30719
rect 14553 30679 14611 30685
rect 6730 30608 6736 30660
rect 6788 30648 6794 30660
rect 7745 30651 7803 30657
rect 7745 30648 7757 30651
rect 6788 30620 7757 30648
rect 6788 30608 6794 30620
rect 7745 30617 7757 30620
rect 7791 30617 7803 30651
rect 7745 30611 7803 30617
rect 9674 30608 9680 30660
rect 9732 30648 9738 30660
rect 14274 30648 14280 30660
rect 9732 30620 14280 30648
rect 9732 30608 9738 30620
rect 14274 30608 14280 30620
rect 14332 30648 14338 30660
rect 14384 30648 14412 30679
rect 14332 30620 14412 30648
rect 14332 30608 14338 30620
rect 7926 30540 7932 30592
rect 7984 30589 7990 30592
rect 7984 30583 8003 30589
rect 7991 30549 8003 30583
rect 7984 30543 8003 30549
rect 7984 30540 7990 30543
rect 10226 30540 10232 30592
rect 10284 30580 10290 30592
rect 14476 30580 14504 30679
rect 14568 30648 14596 30679
rect 14642 30676 14648 30728
rect 14700 30716 14706 30728
rect 14737 30719 14795 30725
rect 14737 30716 14749 30719
rect 14700 30688 14749 30716
rect 14700 30676 14706 30688
rect 14737 30685 14749 30688
rect 14783 30685 14795 30719
rect 14844 30716 14872 30756
rect 15194 30744 15200 30796
rect 15252 30784 15258 30796
rect 15473 30787 15531 30793
rect 15473 30784 15485 30787
rect 15252 30756 15485 30784
rect 15252 30744 15258 30756
rect 15473 30753 15485 30756
rect 15519 30753 15531 30787
rect 17310 30784 17316 30796
rect 17271 30756 17316 30784
rect 15473 30747 15531 30753
rect 17310 30744 17316 30756
rect 17368 30744 17374 30796
rect 19306 30784 19334 30824
rect 19518 30812 19524 30864
rect 19576 30852 19582 30864
rect 19978 30852 19984 30864
rect 19576 30824 19984 30852
rect 19576 30812 19582 30824
rect 19978 30812 19984 30824
rect 20036 30852 20042 30864
rect 25406 30852 25412 30864
rect 20036 30824 25412 30852
rect 20036 30812 20042 30824
rect 25406 30812 25412 30824
rect 25464 30812 25470 30864
rect 19613 30787 19671 30793
rect 19613 30784 19625 30787
rect 19306 30756 19625 30784
rect 19613 30753 19625 30756
rect 19659 30753 19671 30787
rect 19613 30747 19671 30753
rect 22922 30744 22928 30796
rect 22980 30784 22986 30796
rect 25777 30787 25835 30793
rect 22980 30756 24900 30784
rect 22980 30744 22986 30756
rect 19705 30719 19763 30725
rect 19705 30716 19717 30719
rect 14844 30688 19717 30716
rect 14737 30679 14795 30685
rect 19705 30685 19717 30688
rect 19751 30716 19763 30719
rect 22278 30716 22284 30728
rect 19751 30688 22284 30716
rect 19751 30685 19763 30688
rect 19705 30679 19763 30685
rect 22278 30676 22284 30688
rect 22336 30676 22342 30728
rect 23290 30716 23296 30728
rect 23251 30688 23296 30716
rect 23290 30676 23296 30688
rect 23348 30676 23354 30728
rect 23566 30716 23572 30728
rect 23527 30688 23572 30716
rect 23566 30676 23572 30688
rect 23624 30676 23630 30728
rect 24872 30725 24900 30756
rect 25777 30753 25789 30787
rect 25823 30784 25835 30787
rect 26142 30784 26148 30796
rect 25823 30756 26148 30784
rect 25823 30753 25835 30756
rect 25777 30747 25835 30753
rect 26142 30744 26148 30756
rect 26200 30744 26206 30796
rect 28261 30787 28319 30793
rect 28261 30784 28273 30787
rect 26252 30756 28273 30784
rect 24673 30719 24731 30725
rect 24673 30685 24685 30719
rect 24719 30685 24731 30719
rect 24673 30679 24731 30685
rect 24857 30719 24915 30725
rect 24857 30685 24869 30719
rect 24903 30685 24915 30719
rect 24857 30679 24915 30685
rect 24949 30719 25007 30725
rect 24949 30685 24961 30719
rect 24995 30716 25007 30719
rect 25038 30716 25044 30728
rect 24995 30688 25044 30716
rect 24995 30685 25007 30688
rect 24949 30679 25007 30685
rect 15194 30648 15200 30660
rect 14568 30620 15200 30648
rect 15194 30608 15200 30620
rect 15252 30608 15258 30660
rect 15740 30651 15798 30657
rect 15740 30617 15752 30651
rect 15786 30648 15798 30651
rect 16666 30648 16672 30660
rect 15786 30620 16672 30648
rect 15786 30617 15798 30620
rect 15740 30611 15798 30617
rect 16666 30608 16672 30620
rect 16724 30608 16730 30660
rect 17580 30651 17638 30657
rect 17580 30617 17592 30651
rect 17626 30648 17638 30651
rect 17770 30648 17776 30660
rect 17626 30620 17776 30648
rect 17626 30617 17638 30620
rect 17580 30611 17638 30617
rect 17770 30608 17776 30620
rect 17828 30608 17834 30660
rect 19245 30651 19303 30657
rect 19245 30617 19257 30651
rect 19291 30648 19303 30651
rect 19518 30648 19524 30660
rect 19291 30620 19524 30648
rect 19291 30617 19303 30620
rect 19245 30611 19303 30617
rect 19518 30608 19524 30620
rect 19576 30608 19582 30660
rect 24688 30648 24716 30679
rect 25038 30676 25044 30688
rect 25096 30676 25102 30728
rect 25866 30716 25872 30728
rect 25148 30688 25636 30716
rect 25827 30688 25872 30716
rect 25148 30648 25176 30688
rect 24688 30620 25176 30648
rect 25608 30648 25636 30688
rect 25866 30676 25872 30688
rect 25924 30716 25930 30728
rect 26252 30716 26280 30756
rect 28261 30753 28273 30756
rect 28307 30784 28319 30787
rect 28350 30784 28356 30796
rect 28307 30756 28356 30784
rect 28307 30753 28319 30756
rect 28261 30747 28319 30753
rect 28350 30744 28356 30756
rect 28408 30744 28414 30796
rect 25924 30688 26280 30716
rect 28169 30719 28227 30725
rect 25924 30676 25930 30688
rect 28169 30685 28181 30719
rect 28215 30716 28227 30719
rect 28626 30716 28632 30728
rect 28215 30688 28632 30716
rect 28215 30685 28227 30688
rect 28169 30679 28227 30685
rect 28626 30676 28632 30688
rect 28684 30676 28690 30728
rect 26053 30651 26111 30657
rect 26053 30648 26065 30651
rect 25608 30620 26065 30648
rect 26053 30617 26065 30620
rect 26099 30617 26111 30651
rect 26053 30611 26111 30617
rect 16206 30580 16212 30592
rect 10284 30552 16212 30580
rect 10284 30540 10290 30552
rect 16206 30540 16212 30552
rect 16264 30540 16270 30592
rect 16850 30580 16856 30592
rect 16763 30552 16856 30580
rect 16850 30540 16856 30552
rect 16908 30580 16914 30592
rect 18322 30580 18328 30592
rect 16908 30552 18328 30580
rect 16908 30540 16914 30552
rect 18322 30540 18328 30552
rect 18380 30540 18386 30592
rect 19334 30540 19340 30592
rect 19392 30580 19398 30592
rect 19889 30583 19947 30589
rect 19889 30580 19901 30583
rect 19392 30552 19901 30580
rect 19392 30540 19398 30552
rect 19889 30549 19901 30552
rect 19935 30549 19947 30583
rect 19889 30543 19947 30549
rect 22278 30540 22284 30592
rect 22336 30580 22342 30592
rect 22738 30580 22744 30592
rect 22336 30552 22744 30580
rect 22336 30540 22342 30552
rect 22738 30540 22744 30552
rect 22796 30540 22802 30592
rect 23477 30583 23535 30589
rect 23477 30549 23489 30583
rect 23523 30580 23535 30583
rect 24118 30580 24124 30592
rect 23523 30552 24124 30580
rect 23523 30549 23535 30552
rect 23477 30543 23535 30549
rect 24118 30540 24124 30552
rect 24176 30540 24182 30592
rect 24210 30540 24216 30592
rect 24268 30580 24274 30592
rect 25409 30583 25467 30589
rect 25409 30580 25421 30583
rect 24268 30552 25421 30580
rect 24268 30540 24274 30552
rect 25409 30549 25421 30552
rect 25455 30580 25467 30583
rect 27706 30580 27712 30592
rect 25455 30552 27712 30580
rect 25455 30549 25467 30552
rect 25409 30543 25467 30549
rect 27706 30540 27712 30552
rect 27764 30580 27770 30592
rect 27801 30583 27859 30589
rect 27801 30580 27813 30583
rect 27764 30552 27813 30580
rect 27764 30540 27770 30552
rect 27801 30549 27813 30552
rect 27847 30549 27859 30583
rect 27801 30543 27859 30549
rect 28074 30540 28080 30592
rect 28132 30580 28138 30592
rect 28445 30583 28503 30589
rect 28445 30580 28457 30583
rect 28132 30552 28457 30580
rect 28132 30540 28138 30552
rect 28445 30549 28457 30552
rect 28491 30549 28503 30583
rect 28445 30543 28503 30549
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 7282 30336 7288 30388
rect 7340 30376 7346 30388
rect 8113 30379 8171 30385
rect 8113 30376 8125 30379
rect 7340 30348 8125 30376
rect 7340 30336 7346 30348
rect 8113 30345 8125 30348
rect 8159 30345 8171 30379
rect 8113 30339 8171 30345
rect 12526 30336 12532 30388
rect 12584 30376 12590 30388
rect 13446 30376 13452 30388
rect 12584 30348 13452 30376
rect 12584 30336 12590 30348
rect 13446 30336 13452 30348
rect 13504 30336 13510 30388
rect 16206 30336 16212 30388
rect 16264 30376 16270 30388
rect 17218 30376 17224 30388
rect 16264 30348 17224 30376
rect 16264 30336 16270 30348
rect 6362 30268 6368 30320
rect 6420 30308 6426 30320
rect 6730 30308 6736 30320
rect 6420 30280 6736 30308
rect 6420 30268 6426 30280
rect 6730 30268 6736 30280
rect 6788 30308 6794 30320
rect 7745 30311 7803 30317
rect 7745 30308 7757 30311
rect 6788 30280 7757 30308
rect 6788 30268 6794 30280
rect 7745 30277 7757 30280
rect 7791 30277 7803 30311
rect 7926 30308 7932 30320
rect 7984 30317 7990 30320
rect 7984 30311 8019 30317
rect 7871 30280 7932 30308
rect 7745 30271 7803 30277
rect 7926 30268 7932 30280
rect 8007 30308 8019 30311
rect 10870 30308 10876 30320
rect 8007 30280 10876 30308
rect 8007 30277 8019 30280
rect 7984 30271 8019 30277
rect 7984 30268 7990 30271
rect 10870 30268 10876 30280
rect 10928 30268 10934 30320
rect 13630 30308 13636 30320
rect 13591 30280 13636 30308
rect 13630 30268 13636 30280
rect 13688 30268 13694 30320
rect 13814 30268 13820 30320
rect 13872 30308 13878 30320
rect 14642 30308 14648 30320
rect 13872 30280 14648 30308
rect 13872 30268 13878 30280
rect 14642 30268 14648 30280
rect 14700 30268 14706 30320
rect 15194 30308 15200 30320
rect 15155 30280 15200 30308
rect 15194 30268 15200 30280
rect 15252 30268 15258 30320
rect 16666 30308 16672 30320
rect 16627 30280 16672 30308
rect 16666 30268 16672 30280
rect 16724 30268 16730 30320
rect 10502 30200 10508 30252
rect 10560 30240 10566 30252
rect 13449 30243 13507 30249
rect 13449 30240 13461 30243
rect 10560 30212 13461 30240
rect 10560 30200 10566 30212
rect 13449 30209 13461 30212
rect 13495 30209 13507 30243
rect 13449 30203 13507 30209
rect 14829 30243 14887 30249
rect 14829 30209 14841 30243
rect 14875 30209 14887 30243
rect 14829 30203 14887 30209
rect 15013 30243 15071 30249
rect 15013 30209 15025 30243
rect 15059 30240 15071 30243
rect 15654 30240 15660 30252
rect 15059 30212 15660 30240
rect 15059 30209 15071 30212
rect 15013 30203 15071 30209
rect 14844 30172 14872 30203
rect 15654 30200 15660 30212
rect 15712 30240 15718 30252
rect 16942 30240 16948 30252
rect 15712 30212 16620 30240
rect 16903 30212 16948 30240
rect 15712 30200 15718 30212
rect 16482 30172 16488 30184
rect 14844 30144 16488 30172
rect 16482 30132 16488 30144
rect 16540 30132 16546 30184
rect 16592 30172 16620 30212
rect 16942 30200 16948 30212
rect 17000 30200 17006 30252
rect 17052 30249 17080 30348
rect 17218 30336 17224 30348
rect 17276 30336 17282 30388
rect 17770 30376 17776 30388
rect 17731 30348 17776 30376
rect 17770 30336 17776 30348
rect 17828 30336 17834 30388
rect 18506 30376 18512 30388
rect 17880 30348 18512 30376
rect 17037 30243 17095 30249
rect 17037 30209 17049 30243
rect 17083 30209 17095 30243
rect 17037 30203 17095 30209
rect 17126 30200 17132 30252
rect 17184 30240 17190 30252
rect 17184 30212 17229 30240
rect 17184 30200 17190 30212
rect 17310 30200 17316 30252
rect 17368 30240 17374 30252
rect 17368 30212 17413 30240
rect 17368 30200 17374 30212
rect 17880 30172 17908 30348
rect 18506 30336 18512 30348
rect 18564 30336 18570 30388
rect 18782 30376 18788 30388
rect 18743 30348 18788 30376
rect 18782 30336 18788 30348
rect 18840 30336 18846 30388
rect 20806 30336 20812 30388
rect 20864 30376 20870 30388
rect 21634 30376 21640 30388
rect 20864 30348 21640 30376
rect 20864 30336 20870 30348
rect 21634 30336 21640 30348
rect 21692 30336 21698 30388
rect 22094 30336 22100 30388
rect 22152 30376 22158 30388
rect 22649 30379 22707 30385
rect 22649 30376 22661 30379
rect 22152 30348 22661 30376
rect 22152 30336 22158 30348
rect 22649 30345 22661 30348
rect 22695 30376 22707 30379
rect 23566 30376 23572 30388
rect 22695 30348 23572 30376
rect 22695 30345 22707 30348
rect 22649 30339 22707 30345
rect 23566 30336 23572 30348
rect 23624 30336 23630 30388
rect 24581 30379 24639 30385
rect 24581 30345 24593 30379
rect 24627 30376 24639 30379
rect 24946 30376 24952 30388
rect 24627 30348 24952 30376
rect 24627 30345 24639 30348
rect 24581 30339 24639 30345
rect 24946 30336 24952 30348
rect 25004 30376 25010 30388
rect 25130 30376 25136 30388
rect 25004 30348 25136 30376
rect 25004 30336 25010 30348
rect 25130 30336 25136 30348
rect 25188 30336 25194 30388
rect 27798 30336 27804 30388
rect 27856 30376 27862 30388
rect 28261 30379 28319 30385
rect 28261 30376 28273 30379
rect 27856 30348 28273 30376
rect 27856 30336 27862 30348
rect 28261 30345 28273 30348
rect 28307 30376 28319 30379
rect 28810 30376 28816 30388
rect 28307 30348 28816 30376
rect 28307 30345 28319 30348
rect 28261 30339 28319 30345
rect 28810 30336 28816 30348
rect 28868 30336 28874 30388
rect 19334 30308 19340 30320
rect 17972 30280 19340 30308
rect 17972 30249 18000 30280
rect 19334 30268 19340 30280
rect 19392 30268 19398 30320
rect 20625 30311 20683 30317
rect 20625 30277 20637 30311
rect 20671 30308 20683 30311
rect 21818 30308 21824 30320
rect 20671 30280 21824 30308
rect 20671 30277 20683 30280
rect 20625 30271 20683 30277
rect 21818 30268 21824 30280
rect 21876 30268 21882 30320
rect 24486 30308 24492 30320
rect 23032 30280 24492 30308
rect 17957 30243 18015 30249
rect 17957 30209 17969 30243
rect 18003 30209 18015 30243
rect 17957 30203 18015 30209
rect 18141 30243 18199 30249
rect 18141 30209 18153 30243
rect 18187 30209 18199 30243
rect 18141 30203 18199 30209
rect 16592 30144 17908 30172
rect 8570 30104 8576 30116
rect 7944 30076 8576 30104
rect 7944 30045 7972 30076
rect 8570 30064 8576 30076
rect 8628 30064 8634 30116
rect 7929 30039 7987 30045
rect 7929 30005 7941 30039
rect 7975 30005 7987 30039
rect 7929 29999 7987 30005
rect 12986 29996 12992 30048
rect 13044 30036 13050 30048
rect 13630 30036 13636 30048
rect 13044 30008 13636 30036
rect 13044 29996 13050 30008
rect 13630 29996 13636 30008
rect 13688 29996 13694 30048
rect 16298 29996 16304 30048
rect 16356 30036 16362 30048
rect 16942 30036 16948 30048
rect 16356 30008 16948 30036
rect 16356 29996 16362 30008
rect 16942 29996 16948 30008
rect 17000 29996 17006 30048
rect 18156 30036 18184 30203
rect 18230 30200 18236 30252
rect 18288 30240 18294 30252
rect 18288 30212 18333 30240
rect 18288 30200 18294 30212
rect 18506 30200 18512 30252
rect 18564 30240 18570 30252
rect 18693 30243 18751 30249
rect 18693 30240 18705 30243
rect 18564 30212 18705 30240
rect 18564 30200 18570 30212
rect 18693 30209 18705 30212
rect 18739 30209 18751 30243
rect 18693 30203 18751 30209
rect 18877 30243 18935 30249
rect 18877 30209 18889 30243
rect 18923 30209 18935 30243
rect 18877 30203 18935 30209
rect 18322 30132 18328 30184
rect 18380 30172 18386 30184
rect 18892 30172 18920 30203
rect 20346 30200 20352 30252
rect 20404 30240 20410 30252
rect 20441 30243 20499 30249
rect 20441 30240 20453 30243
rect 20404 30212 20453 30240
rect 20404 30200 20410 30212
rect 20441 30209 20453 30212
rect 20487 30209 20499 30243
rect 20441 30203 20499 30209
rect 22557 30243 22615 30249
rect 22557 30209 22569 30243
rect 22603 30240 22615 30243
rect 23032 30240 23060 30280
rect 24486 30268 24492 30280
rect 24544 30308 24550 30320
rect 25961 30311 26019 30317
rect 25961 30308 25973 30311
rect 24544 30280 25973 30308
rect 24544 30268 24550 30280
rect 25961 30277 25973 30280
rect 26007 30277 26019 30311
rect 25961 30271 26019 30277
rect 27893 30311 27951 30317
rect 27893 30277 27905 30311
rect 27939 30308 27951 30311
rect 29178 30308 29184 30320
rect 27939 30280 29184 30308
rect 27939 30277 27951 30280
rect 27893 30271 27951 30277
rect 29178 30268 29184 30280
rect 29236 30268 29242 30320
rect 22603 30212 23060 30240
rect 22603 30209 22615 30212
rect 22557 30203 22615 30209
rect 23106 30200 23112 30252
rect 23164 30240 23170 30252
rect 23457 30243 23515 30249
rect 23457 30240 23469 30243
rect 23164 30212 23469 30240
rect 23164 30200 23170 30212
rect 23457 30209 23469 30212
rect 23503 30209 23515 30243
rect 28074 30240 28080 30252
rect 28035 30212 28080 30240
rect 23457 30203 23515 30209
rect 28074 30200 28080 30212
rect 28132 30200 28138 30252
rect 28337 30233 28395 30239
rect 28337 30230 28349 30233
rect 28276 30202 28349 30230
rect 18380 30144 18920 30172
rect 18380 30132 18386 30144
rect 22186 30132 22192 30184
rect 22244 30172 22250 30184
rect 23201 30175 23259 30181
rect 23201 30172 23213 30175
rect 22244 30144 23213 30172
rect 22244 30132 22250 30144
rect 23201 30141 23213 30144
rect 23247 30141 23259 30175
rect 28276 30172 28304 30202
rect 28337 30199 28349 30202
rect 28383 30199 28395 30233
rect 28337 30193 28395 30199
rect 23201 30135 23259 30141
rect 28092 30144 28304 30172
rect 28092 30116 28120 30144
rect 25866 30104 25872 30116
rect 24504 30076 25872 30104
rect 18322 30036 18328 30048
rect 18156 30008 18328 30036
rect 18322 29996 18328 30008
rect 18380 30036 18386 30048
rect 19426 30036 19432 30048
rect 18380 30008 19432 30036
rect 18380 29996 18386 30008
rect 19426 29996 19432 30008
rect 19484 29996 19490 30048
rect 19518 29996 19524 30048
rect 19576 30036 19582 30048
rect 24504 30036 24532 30076
rect 25866 30064 25872 30076
rect 25924 30064 25930 30116
rect 28074 30064 28080 30116
rect 28132 30064 28138 30116
rect 19576 30008 24532 30036
rect 19576 29996 19582 30008
rect 25774 29996 25780 30048
rect 25832 30036 25838 30048
rect 26053 30039 26111 30045
rect 26053 30036 26065 30039
rect 25832 30008 26065 30036
rect 25832 29996 25838 30008
rect 26053 30005 26065 30008
rect 26099 30005 26111 30039
rect 26053 29999 26111 30005
rect 28258 29996 28264 30048
rect 28316 30036 28322 30048
rect 28902 30036 28908 30048
rect 28316 30008 28908 30036
rect 28316 29996 28322 30008
rect 28902 29996 28908 30008
rect 28960 29996 28966 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 5629 29835 5687 29841
rect 5629 29801 5641 29835
rect 5675 29832 5687 29835
rect 5810 29832 5816 29844
rect 5675 29804 5816 29832
rect 5675 29801 5687 29804
rect 5629 29795 5687 29801
rect 5810 29792 5816 29804
rect 5868 29792 5874 29844
rect 9493 29835 9551 29841
rect 9493 29801 9505 29835
rect 9539 29832 9551 29835
rect 10410 29832 10416 29844
rect 9539 29804 10416 29832
rect 9539 29801 9551 29804
rect 9493 29795 9551 29801
rect 10410 29792 10416 29804
rect 10468 29792 10474 29844
rect 11517 29835 11575 29841
rect 11517 29801 11529 29835
rect 11563 29832 11575 29835
rect 11790 29832 11796 29844
rect 11563 29804 11796 29832
rect 11563 29801 11575 29804
rect 11517 29795 11575 29801
rect 11790 29792 11796 29804
rect 11848 29832 11854 29844
rect 12434 29832 12440 29844
rect 11848 29804 12440 29832
rect 11848 29792 11854 29804
rect 12434 29792 12440 29804
rect 12492 29792 12498 29844
rect 15746 29792 15752 29844
rect 15804 29832 15810 29844
rect 18601 29835 18659 29841
rect 18601 29832 18613 29835
rect 15804 29804 18613 29832
rect 15804 29792 15810 29804
rect 18601 29801 18613 29804
rect 18647 29801 18659 29835
rect 18601 29795 18659 29801
rect 22097 29835 22155 29841
rect 22097 29801 22109 29835
rect 22143 29832 22155 29835
rect 22186 29832 22192 29844
rect 22143 29804 22192 29832
rect 22143 29801 22155 29804
rect 22097 29795 22155 29801
rect 22186 29792 22192 29804
rect 22244 29792 22250 29844
rect 23106 29832 23112 29844
rect 23067 29804 23112 29832
rect 23106 29792 23112 29804
rect 23164 29792 23170 29844
rect 24578 29792 24584 29844
rect 24636 29832 24642 29844
rect 26789 29835 26847 29841
rect 26789 29832 26801 29835
rect 24636 29804 26801 29832
rect 24636 29792 24642 29804
rect 26789 29801 26801 29804
rect 26835 29801 26847 29835
rect 28902 29832 28908 29844
rect 28815 29804 28908 29832
rect 26789 29795 26847 29801
rect 28902 29792 28908 29804
rect 28960 29832 28966 29844
rect 29546 29832 29552 29844
rect 28960 29804 29552 29832
rect 28960 29792 28966 29804
rect 29546 29792 29552 29804
rect 29604 29792 29610 29844
rect 30742 29792 30748 29844
rect 30800 29832 30806 29844
rect 33321 29835 33379 29841
rect 33321 29832 33333 29835
rect 30800 29804 33333 29832
rect 30800 29792 30806 29804
rect 33321 29801 33333 29804
rect 33367 29801 33379 29835
rect 33321 29795 33379 29801
rect 19518 29764 19524 29776
rect 11164 29736 19524 29764
rect 9306 29656 9312 29708
rect 9364 29696 9370 29708
rect 9766 29696 9772 29708
rect 9364 29668 9772 29696
rect 9364 29656 9370 29668
rect 9766 29656 9772 29668
rect 9824 29656 9830 29708
rect 4985 29631 5043 29637
rect 4985 29597 4997 29631
rect 5031 29597 5043 29631
rect 4985 29591 5043 29597
rect 6457 29631 6515 29637
rect 6457 29597 6469 29631
rect 6503 29628 6515 29631
rect 6730 29628 6736 29640
rect 6503 29600 6736 29628
rect 6503 29597 6515 29600
rect 6457 29591 6515 29597
rect 4798 29492 4804 29504
rect 4759 29464 4804 29492
rect 4798 29452 4804 29464
rect 4856 29452 4862 29504
rect 5000 29492 5028 29591
rect 6730 29588 6736 29600
rect 6788 29588 6794 29640
rect 7929 29631 7987 29637
rect 7929 29597 7941 29631
rect 7975 29628 7987 29631
rect 8110 29628 8116 29640
rect 7975 29600 8116 29628
rect 7975 29597 7987 29600
rect 7929 29591 7987 29597
rect 8110 29588 8116 29600
rect 8168 29588 8174 29640
rect 9030 29588 9036 29640
rect 9088 29628 9094 29640
rect 10137 29631 10195 29637
rect 10137 29628 10149 29631
rect 9088 29600 10149 29628
rect 9088 29588 9094 29600
rect 10137 29597 10149 29600
rect 10183 29597 10195 29631
rect 10137 29591 10195 29597
rect 10870 29588 10876 29640
rect 10928 29628 10934 29640
rect 11164 29628 11192 29736
rect 19518 29724 19524 29736
rect 19576 29724 19582 29776
rect 22738 29724 22744 29776
rect 22796 29764 22802 29776
rect 24762 29764 24768 29776
rect 22796 29736 24768 29764
rect 22796 29724 22802 29736
rect 24762 29724 24768 29736
rect 24820 29724 24826 29776
rect 31294 29724 31300 29776
rect 31352 29764 31358 29776
rect 31481 29767 31539 29773
rect 31481 29764 31493 29767
rect 31352 29736 31493 29764
rect 31352 29724 31358 29736
rect 31481 29733 31493 29736
rect 31527 29733 31539 29767
rect 31481 29727 31539 29733
rect 13078 29656 13084 29708
rect 13136 29696 13142 29708
rect 13446 29696 13452 29708
rect 13136 29668 13452 29696
rect 13136 29656 13142 29668
rect 13446 29656 13452 29668
rect 13504 29656 13510 29708
rect 14918 29656 14924 29708
rect 14976 29696 14982 29708
rect 24302 29696 24308 29708
rect 14976 29668 24308 29696
rect 14976 29656 14982 29668
rect 10928 29600 11192 29628
rect 11977 29631 12035 29637
rect 10928 29588 10934 29600
rect 11977 29597 11989 29631
rect 12023 29628 12035 29631
rect 12805 29631 12863 29637
rect 12805 29628 12817 29631
rect 12023 29600 12817 29628
rect 12023 29597 12035 29600
rect 11977 29591 12035 29597
rect 12805 29597 12817 29600
rect 12851 29628 12863 29631
rect 13538 29628 13544 29640
rect 12851 29600 13544 29628
rect 12851 29597 12863 29600
rect 12805 29591 12863 29597
rect 13538 29588 13544 29600
rect 13596 29628 13602 29640
rect 14274 29628 14280 29640
rect 13596 29600 14136 29628
rect 14235 29600 14280 29628
rect 13596 29588 13602 29600
rect 5445 29563 5503 29569
rect 5445 29529 5457 29563
rect 5491 29560 5503 29563
rect 5534 29560 5540 29572
rect 5491 29532 5540 29560
rect 5491 29529 5503 29532
rect 5445 29523 5503 29529
rect 5534 29520 5540 29532
rect 5592 29520 5598 29572
rect 5661 29563 5719 29569
rect 5661 29529 5673 29563
rect 5707 29560 5719 29563
rect 5707 29532 9260 29560
rect 5707 29529 5719 29532
rect 5661 29523 5719 29529
rect 5813 29495 5871 29501
rect 5813 29492 5825 29495
rect 5000 29464 5825 29492
rect 5813 29461 5825 29464
rect 5859 29461 5871 29495
rect 5813 29455 5871 29461
rect 5902 29452 5908 29504
rect 5960 29492 5966 29504
rect 6273 29495 6331 29501
rect 6273 29492 6285 29495
rect 5960 29464 6285 29492
rect 5960 29452 5966 29464
rect 6273 29461 6285 29464
rect 6319 29461 6331 29495
rect 6273 29455 6331 29461
rect 7558 29452 7564 29504
rect 7616 29492 7622 29504
rect 7745 29495 7803 29501
rect 7745 29492 7757 29495
rect 7616 29464 7757 29492
rect 7616 29452 7622 29464
rect 7745 29461 7757 29464
rect 7791 29461 7803 29495
rect 9232 29492 9260 29532
rect 9306 29520 9312 29572
rect 9364 29560 9370 29572
rect 10226 29560 10232 29572
rect 9364 29532 9409 29560
rect 9600 29532 10232 29560
rect 9364 29520 9370 29532
rect 9509 29495 9567 29501
rect 9509 29492 9521 29495
rect 9232 29464 9521 29492
rect 7745 29455 7803 29461
rect 9509 29461 9521 29464
rect 9555 29492 9567 29495
rect 9600 29492 9628 29532
rect 10226 29520 10232 29532
rect 10284 29520 10290 29572
rect 10404 29563 10462 29569
rect 10404 29529 10416 29563
rect 10450 29560 10462 29563
rect 11606 29560 11612 29572
rect 10450 29532 11612 29560
rect 10450 29529 10462 29532
rect 10404 29523 10462 29529
rect 11606 29520 11612 29532
rect 11664 29520 11670 29572
rect 11882 29520 11888 29572
rect 11940 29560 11946 29572
rect 12161 29563 12219 29569
rect 12161 29560 12173 29563
rect 11940 29532 12173 29560
rect 11940 29520 11946 29532
rect 12161 29529 12173 29532
rect 12207 29529 12219 29563
rect 12161 29523 12219 29529
rect 12989 29563 13047 29569
rect 12989 29529 13001 29563
rect 13035 29560 13047 29563
rect 13630 29560 13636 29572
rect 13035 29532 13636 29560
rect 13035 29529 13047 29532
rect 12989 29523 13047 29529
rect 13630 29520 13636 29532
rect 13688 29520 13694 29572
rect 14108 29569 14136 29600
rect 14274 29588 14280 29600
rect 14332 29588 14338 29640
rect 14642 29588 14648 29640
rect 14700 29628 14706 29640
rect 17310 29628 17316 29640
rect 14700 29600 17316 29628
rect 14700 29588 14706 29600
rect 17310 29588 17316 29600
rect 17368 29588 17374 29640
rect 22462 29628 22468 29640
rect 17420 29600 22468 29628
rect 14093 29563 14151 29569
rect 14093 29529 14105 29563
rect 14139 29560 14151 29563
rect 17420 29560 17448 29600
rect 22462 29588 22468 29600
rect 22520 29588 22526 29640
rect 23290 29588 23296 29640
rect 23348 29637 23354 29640
rect 23472 29637 23500 29668
rect 24302 29656 24308 29668
rect 24360 29656 24366 29708
rect 27522 29696 27528 29708
rect 27483 29668 27528 29696
rect 27522 29656 27528 29668
rect 27580 29656 27586 29708
rect 23348 29631 23397 29637
rect 23348 29597 23351 29631
rect 23385 29597 23397 29631
rect 23348 29591 23397 29597
rect 23458 29631 23516 29637
rect 23458 29597 23470 29631
rect 23504 29597 23516 29631
rect 23458 29591 23516 29597
rect 23348 29588 23354 29591
rect 23566 29588 23572 29640
rect 23624 29628 23630 29640
rect 23624 29600 23669 29628
rect 23624 29588 23630 29600
rect 23750 29588 23756 29640
rect 23808 29628 23814 29640
rect 23808 29600 23853 29628
rect 23808 29588 23814 29600
rect 24210 29588 24216 29640
rect 24268 29628 24274 29640
rect 24397 29631 24455 29637
rect 24397 29628 24409 29631
rect 24268 29600 24409 29628
rect 24268 29588 24274 29600
rect 24397 29597 24409 29600
rect 24443 29628 24455 29631
rect 24670 29628 24676 29640
rect 24443 29600 24676 29628
rect 24443 29597 24455 29600
rect 24397 29591 24455 29597
rect 24670 29588 24676 29600
rect 24728 29588 24734 29640
rect 25038 29588 25044 29640
rect 25096 29628 25102 29640
rect 25409 29631 25467 29637
rect 25409 29628 25421 29631
rect 25096 29600 25421 29628
rect 25096 29588 25102 29600
rect 25409 29597 25421 29600
rect 25455 29628 25467 29631
rect 27540 29628 27568 29656
rect 30098 29628 30104 29640
rect 25455 29600 27568 29628
rect 30059 29600 30104 29628
rect 25455 29597 25467 29600
rect 25409 29591 25467 29597
rect 30098 29588 30104 29600
rect 30156 29628 30162 29640
rect 31938 29628 31944 29640
rect 30156 29600 31944 29628
rect 30156 29588 30162 29600
rect 31938 29588 31944 29600
rect 31996 29588 32002 29640
rect 18506 29560 18512 29572
rect 14139 29532 17448 29560
rect 18467 29532 18512 29560
rect 14139 29529 14151 29532
rect 14093 29523 14151 29529
rect 18506 29520 18512 29532
rect 18564 29520 18570 29572
rect 19242 29560 19248 29572
rect 19203 29532 19248 29560
rect 19242 29520 19248 29532
rect 19300 29520 19306 29572
rect 19334 29520 19340 29572
rect 19392 29560 19398 29572
rect 19429 29563 19487 29569
rect 19429 29560 19441 29563
rect 19392 29532 19441 29560
rect 19392 29520 19398 29532
rect 19429 29529 19441 29532
rect 19475 29560 19487 29563
rect 20254 29560 20260 29572
rect 19475 29532 20260 29560
rect 19475 29529 19487 29532
rect 19429 29523 19487 29529
rect 20254 29520 20260 29532
rect 20312 29520 20318 29572
rect 20625 29563 20683 29569
rect 20625 29529 20637 29563
rect 20671 29560 20683 29563
rect 22738 29560 22744 29572
rect 20671 29532 22744 29560
rect 20671 29529 20683 29532
rect 20625 29523 20683 29529
rect 22738 29520 22744 29532
rect 22796 29520 22802 29572
rect 25682 29569 25688 29572
rect 25676 29523 25688 29569
rect 25740 29560 25746 29572
rect 27798 29569 27804 29572
rect 25740 29532 25776 29560
rect 25682 29520 25688 29523
rect 25740 29520 25746 29532
rect 27792 29523 27804 29569
rect 27856 29560 27862 29572
rect 27856 29532 27892 29560
rect 27798 29520 27804 29523
rect 27856 29520 27862 29532
rect 29638 29520 29644 29572
rect 29696 29560 29702 29572
rect 30346 29563 30404 29569
rect 30346 29560 30358 29563
rect 29696 29532 30358 29560
rect 29696 29520 29702 29532
rect 30346 29529 30358 29532
rect 30392 29529 30404 29563
rect 30346 29523 30404 29529
rect 30558 29520 30564 29572
rect 30616 29560 30622 29572
rect 32186 29563 32244 29569
rect 32186 29560 32198 29563
rect 30616 29532 32198 29560
rect 30616 29520 30622 29532
rect 32186 29529 32198 29532
rect 32232 29529 32244 29563
rect 32186 29523 32244 29529
rect 9555 29464 9628 29492
rect 9677 29495 9735 29501
rect 9555 29461 9567 29464
rect 9509 29455 9567 29461
rect 9677 29461 9689 29495
rect 9723 29492 9735 29495
rect 10594 29492 10600 29504
rect 9723 29464 10600 29492
rect 9723 29461 9735 29464
rect 9677 29455 9735 29461
rect 10594 29452 10600 29464
rect 10652 29452 10658 29504
rect 12066 29452 12072 29504
rect 12124 29492 12130 29504
rect 12345 29495 12403 29501
rect 12345 29492 12357 29495
rect 12124 29464 12357 29492
rect 12124 29452 12130 29464
rect 12345 29461 12357 29464
rect 12391 29461 12403 29495
rect 13170 29492 13176 29504
rect 13131 29464 13176 29492
rect 12345 29455 12403 29461
rect 13170 29452 13176 29464
rect 13228 29452 13234 29504
rect 14461 29495 14519 29501
rect 14461 29461 14473 29495
rect 14507 29492 14519 29495
rect 14826 29492 14832 29504
rect 14507 29464 14832 29492
rect 14507 29461 14519 29464
rect 14461 29455 14519 29461
rect 14826 29452 14832 29464
rect 14884 29452 14890 29504
rect 19613 29495 19671 29501
rect 19613 29461 19625 29495
rect 19659 29492 19671 29495
rect 21174 29492 21180 29504
rect 19659 29464 21180 29492
rect 19659 29461 19671 29464
rect 19613 29455 19671 29461
rect 21174 29452 21180 29464
rect 21232 29452 21238 29504
rect 23750 29452 23756 29504
rect 23808 29492 23814 29504
rect 24581 29495 24639 29501
rect 24581 29492 24593 29495
rect 23808 29464 24593 29492
rect 23808 29452 23814 29464
rect 24581 29461 24593 29464
rect 24627 29461 24639 29495
rect 24581 29455 24639 29461
rect 24670 29452 24676 29504
rect 24728 29492 24734 29504
rect 26970 29492 26976 29504
rect 24728 29464 26976 29492
rect 24728 29452 24734 29464
rect 26970 29452 26976 29464
rect 27028 29452 27034 29504
rect 30466 29452 30472 29504
rect 30524 29492 30530 29504
rect 31294 29492 31300 29504
rect 30524 29464 31300 29492
rect 30524 29452 30530 29464
rect 31294 29452 31300 29464
rect 31352 29452 31358 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 5534 29288 5540 29300
rect 4632 29260 5540 29288
rect 4433 29155 4491 29161
rect 4433 29121 4445 29155
rect 4479 29152 4491 29155
rect 4632 29152 4660 29260
rect 5534 29248 5540 29260
rect 5592 29288 5598 29300
rect 6822 29288 6828 29300
rect 5592 29260 6828 29288
rect 5592 29248 5598 29260
rect 6822 29248 6828 29260
rect 6880 29248 6886 29300
rect 10410 29288 10416 29300
rect 10371 29260 10416 29288
rect 10410 29248 10416 29260
rect 10468 29248 10474 29300
rect 11606 29288 11612 29300
rect 11567 29260 11612 29288
rect 11606 29248 11612 29260
rect 11664 29248 11670 29300
rect 11882 29248 11888 29300
rect 11940 29288 11946 29300
rect 13078 29288 13084 29300
rect 11940 29260 13084 29288
rect 11940 29248 11946 29260
rect 13078 29248 13084 29260
rect 13136 29248 13142 29300
rect 14090 29288 14096 29300
rect 14051 29260 14096 29288
rect 14090 29248 14096 29260
rect 14148 29248 14154 29300
rect 15838 29248 15844 29300
rect 15896 29288 15902 29300
rect 15933 29291 15991 29297
rect 15933 29288 15945 29291
rect 15896 29260 15945 29288
rect 15896 29248 15902 29260
rect 15933 29257 15945 29260
rect 15979 29257 15991 29291
rect 15933 29251 15991 29257
rect 22002 29248 22008 29300
rect 22060 29288 22066 29300
rect 22830 29288 22836 29300
rect 22060 29260 22836 29288
rect 22060 29248 22066 29260
rect 22830 29248 22836 29260
rect 22888 29288 22894 29300
rect 23201 29291 23259 29297
rect 23201 29288 23213 29291
rect 22888 29260 23213 29288
rect 22888 29248 22894 29260
rect 23201 29257 23213 29260
rect 23247 29257 23259 29291
rect 23201 29251 23259 29257
rect 23566 29248 23572 29300
rect 23624 29288 23630 29300
rect 24029 29291 24087 29297
rect 24029 29288 24041 29291
rect 23624 29260 24041 29288
rect 23624 29248 23630 29260
rect 24029 29257 24041 29260
rect 24075 29257 24087 29291
rect 24029 29251 24087 29257
rect 24578 29248 24584 29300
rect 24636 29288 24642 29300
rect 25409 29291 25467 29297
rect 24636 29260 25259 29288
rect 24636 29248 24642 29260
rect 4700 29223 4758 29229
rect 4700 29189 4712 29223
rect 4746 29220 4758 29223
rect 4798 29220 4804 29232
rect 4746 29192 4804 29220
rect 4746 29189 4758 29192
rect 4700 29183 4758 29189
rect 4798 29180 4804 29192
rect 4856 29180 4862 29232
rect 6362 29220 6368 29232
rect 6323 29192 6368 29220
rect 6362 29180 6368 29192
rect 6420 29180 6426 29232
rect 6546 29180 6552 29232
rect 6604 29229 6610 29232
rect 6604 29223 6623 29229
rect 6611 29220 6623 29223
rect 7926 29220 7932 29232
rect 6611 29192 7932 29220
rect 6611 29189 6623 29192
rect 6604 29183 6623 29189
rect 6604 29180 6610 29183
rect 7926 29180 7932 29192
rect 7984 29220 7990 29232
rect 10134 29220 10140 29232
rect 7984 29192 8064 29220
rect 7984 29180 7990 29192
rect 8036 29161 8064 29192
rect 9140 29192 10140 29220
rect 4479 29124 4660 29152
rect 8021 29155 8079 29161
rect 4479 29121 4491 29124
rect 4433 29115 4491 29121
rect 8021 29121 8033 29155
rect 8067 29121 8079 29155
rect 9030 29152 9036 29164
rect 8991 29124 9036 29152
rect 8021 29115 8079 29121
rect 9030 29112 9036 29124
rect 9088 29112 9094 29164
rect 7745 29087 7803 29093
rect 7745 29053 7757 29087
rect 7791 29084 7803 29087
rect 9140 29084 9168 29192
rect 10134 29180 10140 29192
rect 10192 29220 10198 29232
rect 10502 29220 10508 29232
rect 10192 29192 10508 29220
rect 10192 29180 10198 29192
rect 10502 29180 10508 29192
rect 10560 29180 10566 29232
rect 12342 29220 12348 29232
rect 11992 29192 12348 29220
rect 9300 29155 9358 29161
rect 9300 29121 9312 29155
rect 9346 29152 9358 29155
rect 10410 29152 10416 29164
rect 9346 29124 10416 29152
rect 9346 29121 9358 29124
rect 9300 29115 9358 29121
rect 10410 29112 10416 29124
rect 10468 29112 10474 29164
rect 11790 29112 11796 29164
rect 11848 29152 11854 29164
rect 11992 29161 12020 29192
rect 12342 29180 12348 29192
rect 12400 29180 12406 29232
rect 12434 29180 12440 29232
rect 12492 29220 12498 29232
rect 12492 29192 14596 29220
rect 12492 29180 12498 29192
rect 11885 29155 11943 29161
rect 11885 29152 11897 29155
rect 11848 29124 11897 29152
rect 11848 29112 11854 29124
rect 11885 29121 11897 29124
rect 11931 29121 11943 29155
rect 11885 29115 11943 29121
rect 11977 29155 12035 29161
rect 11977 29121 11989 29155
rect 12023 29121 12035 29155
rect 11977 29115 12035 29121
rect 12066 29112 12072 29164
rect 12124 29152 12130 29164
rect 12728 29161 12756 29192
rect 12253 29155 12311 29161
rect 12124 29124 12169 29152
rect 12124 29112 12130 29124
rect 12253 29121 12265 29155
rect 12299 29152 12311 29155
rect 12713 29155 12771 29161
rect 12299 29124 12664 29152
rect 12299 29121 12311 29124
rect 12253 29115 12311 29121
rect 7791 29056 9168 29084
rect 7791 29053 7803 29056
rect 7745 29047 7803 29053
rect 5810 29016 5816 29028
rect 5771 28988 5816 29016
rect 5810 28976 5816 28988
rect 5868 28976 5874 29028
rect 6730 29016 6736 29028
rect 6691 28988 6736 29016
rect 6730 28976 6736 28988
rect 6788 28976 6794 29028
rect 6546 28948 6552 28960
rect 6507 28920 6552 28948
rect 6546 28908 6552 28920
rect 6604 28908 6610 28960
rect 11882 28908 11888 28960
rect 11940 28948 11946 28960
rect 12636 28948 12664 29124
rect 12713 29121 12725 29155
rect 12759 29121 12771 29155
rect 12713 29115 12771 29121
rect 12802 29112 12808 29164
rect 12860 29152 12866 29164
rect 14568 29161 14596 29192
rect 15470 29180 15476 29232
rect 15528 29220 15534 29232
rect 15746 29220 15752 29232
rect 15528 29192 15752 29220
rect 15528 29180 15534 29192
rect 15746 29180 15752 29192
rect 15804 29180 15810 29232
rect 20714 29220 20720 29232
rect 19260 29192 20720 29220
rect 12969 29155 13027 29161
rect 12969 29152 12981 29155
rect 12860 29124 12981 29152
rect 12860 29112 12866 29124
rect 12969 29121 12981 29124
rect 13015 29121 13027 29155
rect 12969 29115 13027 29121
rect 14553 29155 14611 29161
rect 14553 29121 14565 29155
rect 14599 29121 14611 29155
rect 14553 29115 14611 29121
rect 14642 29112 14648 29164
rect 14700 29152 14706 29164
rect 14809 29155 14867 29161
rect 14809 29152 14821 29155
rect 14700 29124 14821 29152
rect 14700 29112 14706 29124
rect 14809 29121 14821 29124
rect 14855 29121 14867 29155
rect 14809 29115 14867 29121
rect 17770 29112 17776 29164
rect 17828 29152 17834 29164
rect 19260 29161 19288 29192
rect 20714 29180 20720 29192
rect 20772 29220 20778 29232
rect 21910 29220 21916 29232
rect 20772 29192 21916 29220
rect 20772 29180 20778 29192
rect 17865 29155 17923 29161
rect 17865 29152 17877 29155
rect 17828 29124 17877 29152
rect 17828 29112 17834 29124
rect 17865 29121 17877 29124
rect 17911 29121 17923 29155
rect 17865 29115 17923 29121
rect 19245 29155 19303 29161
rect 19245 29121 19257 29155
rect 19291 29121 19303 29155
rect 19245 29115 19303 29121
rect 19512 29155 19570 29161
rect 19512 29121 19524 29155
rect 19558 29152 19570 29155
rect 20806 29152 20812 29164
rect 19558 29124 20812 29152
rect 19558 29121 19570 29124
rect 19512 29115 19570 29121
rect 20806 29112 20812 29124
rect 20864 29112 20870 29164
rect 21836 29161 21864 29192
rect 21910 29180 21916 29192
rect 21968 29220 21974 29232
rect 22186 29220 22192 29232
rect 21968 29192 22192 29220
rect 21968 29180 21974 29192
rect 22186 29180 22192 29192
rect 22244 29180 22250 29232
rect 24302 29180 24308 29232
rect 24360 29220 24366 29232
rect 24765 29223 24823 29229
rect 24765 29220 24777 29223
rect 24360 29192 24777 29220
rect 24360 29180 24366 29192
rect 24765 29189 24777 29192
rect 24811 29189 24823 29223
rect 24765 29183 24823 29189
rect 22094 29161 22100 29164
rect 21821 29155 21879 29161
rect 21821 29121 21833 29155
rect 21867 29121 21879 29155
rect 21821 29115 21879 29121
rect 22088 29115 22100 29161
rect 22152 29152 22158 29164
rect 22152 29124 22188 29152
rect 22094 29112 22100 29115
rect 22152 29112 22158 29124
rect 22462 29112 22468 29164
rect 22520 29152 22526 29164
rect 23661 29155 23719 29161
rect 23661 29152 23673 29155
rect 22520 29124 23673 29152
rect 22520 29112 22526 29124
rect 23661 29121 23673 29124
rect 23707 29121 23719 29155
rect 23842 29152 23848 29164
rect 23803 29124 23848 29152
rect 23661 29115 23719 29121
rect 17402 29044 17408 29096
rect 17460 29084 17466 29096
rect 17586 29084 17592 29096
rect 17460 29056 17592 29084
rect 17460 29044 17466 29056
rect 17586 29044 17592 29056
rect 17644 29084 17650 29096
rect 17681 29087 17739 29093
rect 17681 29084 17693 29087
rect 17644 29056 17693 29084
rect 17644 29044 17650 29056
rect 17681 29053 17693 29056
rect 17727 29053 17739 29087
rect 23676 29084 23704 29115
rect 23842 29112 23848 29124
rect 23900 29112 23906 29164
rect 24486 29112 24492 29164
rect 24544 29152 24550 29164
rect 24581 29155 24639 29161
rect 24581 29152 24593 29155
rect 24544 29124 24593 29152
rect 24544 29112 24550 29124
rect 24581 29121 24593 29124
rect 24627 29152 24639 29155
rect 24670 29152 24676 29164
rect 24627 29124 24676 29152
rect 24627 29121 24639 29124
rect 24581 29115 24639 29121
rect 24670 29112 24676 29124
rect 24728 29112 24734 29164
rect 25231 29152 25259 29260
rect 25409 29257 25421 29291
rect 25455 29288 25467 29291
rect 25682 29288 25688 29300
rect 25455 29260 25688 29288
rect 25455 29257 25467 29260
rect 25409 29251 25467 29257
rect 25682 29248 25688 29260
rect 25740 29248 25746 29300
rect 27706 29288 27712 29300
rect 27667 29260 27712 29288
rect 27706 29248 27712 29260
rect 27764 29248 27770 29300
rect 29638 29288 29644 29300
rect 29599 29260 29644 29288
rect 29638 29248 29644 29260
rect 29696 29248 29702 29300
rect 30466 29288 30472 29300
rect 30024 29260 30472 29288
rect 30024 29220 30052 29260
rect 30466 29248 30472 29260
rect 30524 29248 30530 29300
rect 25792 29192 29776 29220
rect 25792 29164 25820 29192
rect 25639 29155 25697 29161
rect 25639 29152 25651 29155
rect 25231 29124 25651 29152
rect 25639 29121 25651 29124
rect 25685 29121 25697 29155
rect 25774 29152 25780 29164
rect 25735 29124 25780 29152
rect 25639 29115 25697 29121
rect 25774 29112 25780 29124
rect 25832 29112 25838 29164
rect 25866 29112 25872 29164
rect 25924 29152 25930 29164
rect 26050 29152 26056 29164
rect 25924 29124 25969 29152
rect 26011 29124 26056 29152
rect 25924 29112 25930 29124
rect 26050 29112 26056 29124
rect 26108 29112 26114 29164
rect 28813 29155 28871 29161
rect 28813 29152 28825 29155
rect 26160 29124 28825 29152
rect 26160 29084 26188 29124
rect 28813 29121 28825 29124
rect 28859 29121 28871 29155
rect 28813 29115 28871 29121
rect 28997 29155 29055 29161
rect 28997 29121 29009 29155
rect 29043 29152 29055 29155
rect 29638 29152 29644 29164
rect 29043 29124 29644 29152
rect 29043 29121 29055 29124
rect 28997 29115 29055 29121
rect 29638 29112 29644 29124
rect 29696 29112 29702 29164
rect 23676 29056 26188 29084
rect 28077 29087 28135 29093
rect 17681 29047 17739 29053
rect 28077 29053 28089 29087
rect 28123 29053 28135 29087
rect 28077 29047 28135 29053
rect 28169 29087 28227 29093
rect 28169 29053 28181 29087
rect 28215 29084 28227 29087
rect 28350 29084 28356 29096
rect 28215 29056 28356 29084
rect 28215 29053 28227 29056
rect 28169 29047 28227 29053
rect 18049 29019 18107 29025
rect 18049 28985 18061 29019
rect 18095 29016 18107 29019
rect 18506 29016 18512 29028
rect 18095 28988 18512 29016
rect 18095 28985 18107 28988
rect 18049 28979 18107 28985
rect 18506 28976 18512 28988
rect 18564 29016 18570 29028
rect 18564 28988 19288 29016
rect 18564 28976 18570 28988
rect 14182 28948 14188 28960
rect 11940 28920 14188 28948
rect 11940 28908 11946 28920
rect 14182 28908 14188 28920
rect 14240 28908 14246 28960
rect 15194 28908 15200 28960
rect 15252 28948 15258 28960
rect 15470 28948 15476 28960
rect 15252 28920 15476 28948
rect 15252 28908 15258 28920
rect 15470 28908 15476 28920
rect 15528 28908 15534 28960
rect 19260 28948 19288 28988
rect 20530 28976 20536 29028
rect 20588 29016 20594 29028
rect 20625 29019 20683 29025
rect 20625 29016 20637 29019
rect 20588 28988 20637 29016
rect 20588 28976 20594 28988
rect 20625 28985 20637 28988
rect 20671 29016 20683 29019
rect 21542 29016 21548 29028
rect 20671 28988 21548 29016
rect 20671 28985 20683 28988
rect 20625 28979 20683 28985
rect 21542 28976 21548 28988
rect 21600 28976 21606 29028
rect 23290 28976 23296 29028
rect 23348 29016 23354 29028
rect 25774 29016 25780 29028
rect 23348 28988 25780 29016
rect 23348 28976 23354 28988
rect 25774 28976 25780 28988
rect 25832 28976 25838 29028
rect 25958 28976 25964 29028
rect 26016 28976 26022 29028
rect 28092 29016 28120 29047
rect 28350 29044 28356 29056
rect 28408 29044 28414 29096
rect 29748 29084 29776 29192
rect 29932 29192 30052 29220
rect 29932 29161 29960 29192
rect 29917 29155 29975 29161
rect 29917 29121 29929 29155
rect 29963 29121 29975 29155
rect 29917 29115 29975 29121
rect 30009 29155 30067 29161
rect 30009 29121 30021 29155
rect 30055 29121 30067 29155
rect 30009 29115 30067 29121
rect 30101 29155 30159 29161
rect 30101 29121 30113 29155
rect 30147 29121 30159 29155
rect 30282 29152 30288 29164
rect 30243 29124 30288 29152
rect 30101 29115 30159 29121
rect 29822 29084 29828 29096
rect 29735 29056 29828 29084
rect 29822 29044 29828 29056
rect 29880 29084 29886 29096
rect 30024 29084 30052 29115
rect 29880 29056 30052 29084
rect 30116 29084 30144 29115
rect 30282 29112 30288 29124
rect 30340 29112 30346 29164
rect 31018 29084 31024 29096
rect 30116 29056 31024 29084
rect 29880 29044 29886 29056
rect 31018 29044 31024 29056
rect 31076 29044 31082 29096
rect 28902 29016 28908 29028
rect 28092 28988 28908 29016
rect 28902 28976 28908 28988
rect 28960 28976 28966 29028
rect 29181 29019 29239 29025
rect 29181 28985 29193 29019
rect 29227 29016 29239 29019
rect 30190 29016 30196 29028
rect 29227 28988 30196 29016
rect 29227 28985 29239 28988
rect 29181 28979 29239 28985
rect 30190 28976 30196 28988
rect 30248 28976 30254 29028
rect 30282 28976 30288 29028
rect 30340 28976 30346 29028
rect 19886 28948 19892 28960
rect 19260 28920 19892 28948
rect 19886 28908 19892 28920
rect 19944 28908 19950 28960
rect 22462 28908 22468 28960
rect 22520 28948 22526 28960
rect 25976 28948 26004 28976
rect 27522 28948 27528 28960
rect 22520 28920 27528 28948
rect 22520 28908 22526 28920
rect 27522 28908 27528 28920
rect 27580 28908 27586 28960
rect 27890 28908 27896 28960
rect 27948 28948 27954 28960
rect 28353 28951 28411 28957
rect 28353 28948 28365 28951
rect 27948 28920 28365 28948
rect 27948 28908 27954 28920
rect 28353 28917 28365 28920
rect 28399 28917 28411 28951
rect 28353 28911 28411 28917
rect 29914 28908 29920 28960
rect 29972 28948 29978 28960
rect 30300 28948 30328 28976
rect 29972 28920 30328 28948
rect 29972 28908 29978 28920
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 6822 28744 6828 28756
rect 6783 28716 6828 28744
rect 6822 28704 6828 28716
rect 6880 28704 6886 28756
rect 7929 28747 7987 28753
rect 7929 28713 7941 28747
rect 7975 28744 7987 28747
rect 8662 28744 8668 28756
rect 7975 28716 8668 28744
rect 7975 28713 7987 28716
rect 7929 28707 7987 28713
rect 8662 28704 8668 28716
rect 8720 28704 8726 28756
rect 12713 28747 12771 28753
rect 12713 28713 12725 28747
rect 12759 28744 12771 28747
rect 12802 28744 12808 28756
rect 12759 28716 12808 28744
rect 12759 28713 12771 28716
rect 12713 28707 12771 28713
rect 12802 28704 12808 28716
rect 12860 28704 12866 28756
rect 14553 28747 14611 28753
rect 14553 28713 14565 28747
rect 14599 28744 14611 28747
rect 14642 28744 14648 28756
rect 14599 28716 14648 28744
rect 14599 28713 14611 28716
rect 14553 28707 14611 28713
rect 14642 28704 14648 28716
rect 14700 28704 14706 28756
rect 15010 28744 15016 28756
rect 14752 28716 15016 28744
rect 8110 28676 8116 28688
rect 8071 28648 8116 28676
rect 8110 28636 8116 28648
rect 8168 28636 8174 28688
rect 14090 28608 14096 28620
rect 13004 28580 14096 28608
rect 5537 28543 5595 28549
rect 5537 28509 5549 28543
rect 5583 28540 5595 28543
rect 9490 28540 9496 28552
rect 5583 28512 9496 28540
rect 5583 28509 5595 28512
rect 5537 28503 5595 28509
rect 9490 28500 9496 28512
rect 9548 28540 9554 28552
rect 13004 28549 13032 28580
rect 14090 28568 14096 28580
rect 14148 28568 14154 28620
rect 14752 28608 14780 28716
rect 15010 28704 15016 28716
rect 15068 28704 15074 28756
rect 16114 28744 16120 28756
rect 15304 28716 16120 28744
rect 14826 28636 14832 28688
rect 14884 28676 14890 28688
rect 15304 28676 15332 28716
rect 16114 28704 16120 28716
rect 16172 28744 16178 28756
rect 20438 28744 20444 28756
rect 16172 28716 20444 28744
rect 16172 28704 16178 28716
rect 20438 28704 20444 28716
rect 20496 28704 20502 28756
rect 20717 28747 20775 28753
rect 20717 28713 20729 28747
rect 20763 28744 20775 28747
rect 20806 28744 20812 28756
rect 20763 28716 20812 28744
rect 20763 28713 20775 28716
rect 20717 28707 20775 28713
rect 20806 28704 20812 28716
rect 20864 28704 20870 28756
rect 21821 28747 21879 28753
rect 21821 28713 21833 28747
rect 21867 28744 21879 28747
rect 22094 28744 22100 28756
rect 21867 28716 22100 28744
rect 21867 28713 21879 28716
rect 21821 28707 21879 28713
rect 22094 28704 22100 28716
rect 22152 28704 22158 28756
rect 23290 28744 23296 28756
rect 22195 28716 23296 28744
rect 18046 28676 18052 28688
rect 14884 28648 15056 28676
rect 14884 28636 14890 28648
rect 14752 28580 14955 28608
rect 10505 28543 10563 28549
rect 10505 28540 10517 28543
rect 9548 28512 10517 28540
rect 9548 28500 9554 28512
rect 10505 28509 10517 28512
rect 10551 28509 10563 28543
rect 10505 28503 10563 28509
rect 12989 28543 13047 28549
rect 12989 28509 13001 28543
rect 13035 28509 13047 28543
rect 12989 28503 13047 28509
rect 13081 28543 13139 28549
rect 13081 28509 13093 28543
rect 13127 28509 13139 28543
rect 13081 28503 13139 28509
rect 7742 28472 7748 28484
rect 7703 28444 7748 28472
rect 7742 28432 7748 28444
rect 7800 28432 7806 28484
rect 7926 28432 7932 28484
rect 7984 28481 7990 28484
rect 7984 28475 8003 28481
rect 7991 28441 8003 28475
rect 7984 28435 8003 28441
rect 7984 28432 7990 28435
rect 12710 28432 12716 28484
rect 12768 28472 12774 28484
rect 13096 28472 13124 28503
rect 13170 28500 13176 28552
rect 13228 28540 13234 28552
rect 13357 28543 13415 28549
rect 13228 28512 13273 28540
rect 13228 28500 13234 28512
rect 13357 28509 13369 28543
rect 13403 28540 13415 28543
rect 14182 28540 14188 28552
rect 13403 28512 14188 28540
rect 13403 28509 13415 28512
rect 13357 28503 13415 28509
rect 14182 28500 14188 28512
rect 14240 28500 14246 28552
rect 14752 28472 14780 28580
rect 14927 28549 14955 28580
rect 15028 28549 15056 28648
rect 15212 28648 15332 28676
rect 17144 28648 18052 28676
rect 15212 28549 15240 28648
rect 15470 28568 15476 28620
rect 15528 28608 15534 28620
rect 15749 28611 15807 28617
rect 15749 28608 15761 28611
rect 15528 28580 15761 28608
rect 15528 28568 15534 28580
rect 15749 28577 15761 28580
rect 15795 28577 15807 28611
rect 15749 28571 15807 28577
rect 14829 28543 14887 28549
rect 14829 28509 14841 28543
rect 14875 28509 14887 28543
rect 14829 28503 14887 28509
rect 14918 28543 14976 28549
rect 14918 28509 14930 28543
rect 14964 28509 14976 28543
rect 14918 28503 14976 28509
rect 15018 28543 15076 28549
rect 15018 28509 15030 28543
rect 15064 28509 15076 28543
rect 15018 28503 15076 28509
rect 15197 28543 15255 28549
rect 15197 28509 15209 28543
rect 15243 28509 15255 28543
rect 15838 28540 15844 28552
rect 15197 28503 15255 28509
rect 15396 28512 15844 28540
rect 12768 28444 14780 28472
rect 14844 28472 14872 28503
rect 15396 28472 15424 28512
rect 15838 28500 15844 28512
rect 15896 28500 15902 28552
rect 14844 28444 15424 28472
rect 12768 28432 12774 28444
rect 15470 28432 15476 28484
rect 15528 28472 15534 28484
rect 15994 28475 16052 28481
rect 15994 28472 16006 28475
rect 15528 28444 16006 28472
rect 15528 28432 15534 28444
rect 15994 28441 16006 28444
rect 16040 28441 16052 28475
rect 15994 28435 16052 28441
rect 9030 28364 9036 28416
rect 9088 28404 9094 28416
rect 11514 28404 11520 28416
rect 9088 28376 11520 28404
rect 9088 28364 9094 28376
rect 11514 28364 11520 28376
rect 11572 28404 11578 28416
rect 11793 28407 11851 28413
rect 11793 28404 11805 28407
rect 11572 28376 11805 28404
rect 11572 28364 11578 28376
rect 11793 28373 11805 28376
rect 11839 28404 11851 28407
rect 12158 28404 12164 28416
rect 11839 28376 12164 28404
rect 11839 28373 11851 28376
rect 11793 28367 11851 28373
rect 12158 28364 12164 28376
rect 12216 28364 12222 28416
rect 16758 28364 16764 28416
rect 16816 28404 16822 28416
rect 17144 28413 17172 28648
rect 18046 28636 18052 28648
rect 18104 28636 18110 28688
rect 18601 28679 18659 28685
rect 18601 28645 18613 28679
rect 18647 28676 18659 28679
rect 18647 28648 20392 28676
rect 18647 28645 18659 28648
rect 18601 28639 18659 28645
rect 17954 28568 17960 28620
rect 18012 28608 18018 28620
rect 18012 28580 18460 28608
rect 18012 28568 18018 28580
rect 18046 28540 18052 28552
rect 18007 28512 18052 28540
rect 18046 28500 18052 28512
rect 18104 28500 18110 28552
rect 18432 28549 18460 28580
rect 19794 28568 19800 28620
rect 19852 28608 19858 28620
rect 19852 28580 20024 28608
rect 19852 28568 19858 28580
rect 18417 28543 18475 28549
rect 18417 28509 18429 28543
rect 18463 28509 18475 28543
rect 19518 28540 19524 28552
rect 18417 28503 18475 28509
rect 19306 28512 19524 28540
rect 18230 28472 18236 28484
rect 18191 28444 18236 28472
rect 18230 28432 18236 28444
rect 18288 28432 18294 28484
rect 18325 28475 18383 28481
rect 18325 28441 18337 28475
rect 18371 28472 18383 28475
rect 19306 28472 19334 28512
rect 19518 28500 19524 28512
rect 19576 28500 19582 28552
rect 19702 28540 19708 28552
rect 19663 28512 19708 28540
rect 19702 28500 19708 28512
rect 19760 28500 19766 28552
rect 19886 28540 19892 28552
rect 19847 28512 19892 28540
rect 19886 28500 19892 28512
rect 19944 28500 19950 28552
rect 19996 28549 20024 28580
rect 19981 28543 20039 28549
rect 19981 28509 19993 28543
rect 20027 28509 20039 28543
rect 19981 28503 20039 28509
rect 20165 28543 20223 28549
rect 20165 28509 20177 28543
rect 20211 28509 20223 28543
rect 20165 28503 20223 28509
rect 20257 28543 20315 28549
rect 20257 28509 20269 28543
rect 20303 28540 20315 28543
rect 20364 28540 20392 28648
rect 21542 28636 21548 28688
rect 21600 28676 21606 28688
rect 22002 28676 22008 28688
rect 21600 28648 22008 28676
rect 21600 28636 21606 28648
rect 22002 28636 22008 28648
rect 22060 28636 22066 28688
rect 22195 28608 22223 28716
rect 23290 28704 23296 28716
rect 23348 28704 23354 28756
rect 24581 28747 24639 28753
rect 24581 28713 24593 28747
rect 24627 28713 24639 28747
rect 24581 28707 24639 28713
rect 25685 28747 25743 28753
rect 25685 28713 25697 28747
rect 25731 28744 25743 28747
rect 25866 28744 25872 28756
rect 25731 28716 25872 28744
rect 25731 28713 25743 28716
rect 25685 28707 25743 28713
rect 23293 28611 23351 28617
rect 23293 28608 23305 28611
rect 21100 28580 22232 28608
rect 20303 28512 20392 28540
rect 20303 28509 20315 28512
rect 20257 28503 20315 28509
rect 18371 28444 19334 28472
rect 20180 28472 20208 28503
rect 20530 28500 20536 28552
rect 20588 28540 20594 28552
rect 21100 28549 21128 28580
rect 20993 28543 21051 28549
rect 20993 28540 21005 28543
rect 20588 28512 21005 28540
rect 20588 28500 20594 28512
rect 20993 28509 21005 28512
rect 21039 28509 21051 28543
rect 20993 28503 21051 28509
rect 21085 28543 21143 28549
rect 21085 28509 21097 28543
rect 21131 28509 21143 28543
rect 21085 28503 21143 28509
rect 21174 28500 21180 28552
rect 21232 28540 21238 28552
rect 21361 28543 21419 28549
rect 21232 28512 21277 28540
rect 21232 28500 21238 28512
rect 21361 28509 21373 28543
rect 21407 28509 21419 28543
rect 21361 28503 21419 28509
rect 20898 28472 20904 28484
rect 20180 28444 20904 28472
rect 18371 28441 18383 28444
rect 18325 28435 18383 28441
rect 20898 28432 20904 28444
rect 20956 28432 20962 28484
rect 21376 28472 21404 28503
rect 21542 28500 21548 28552
rect 21600 28540 21606 28552
rect 22204 28549 22232 28580
rect 22296 28580 23305 28608
rect 22296 28549 22324 28580
rect 23293 28577 23305 28580
rect 23339 28577 23351 28611
rect 24596 28608 24624 28707
rect 25866 28704 25872 28716
rect 25924 28704 25930 28756
rect 27617 28747 27675 28753
rect 27617 28713 27629 28747
rect 27663 28744 27675 28747
rect 27798 28744 27804 28756
rect 27663 28716 27804 28744
rect 27663 28713 27675 28716
rect 27617 28707 27675 28713
rect 27798 28704 27804 28716
rect 27856 28704 27862 28756
rect 29733 28747 29791 28753
rect 29733 28713 29745 28747
rect 29779 28744 29791 28747
rect 30558 28744 30564 28756
rect 29779 28716 30564 28744
rect 29779 28713 29791 28716
rect 29733 28707 29791 28713
rect 30558 28704 30564 28716
rect 30616 28704 30622 28756
rect 31938 28704 31944 28756
rect 31996 28744 32002 28756
rect 32401 28747 32459 28753
rect 32401 28744 32413 28747
rect 31996 28716 32413 28744
rect 31996 28704 32002 28716
rect 32401 28713 32413 28716
rect 32447 28713 32459 28747
rect 32401 28707 32459 28713
rect 27522 28636 27528 28688
rect 27580 28676 27586 28688
rect 28813 28679 28871 28685
rect 28813 28676 28825 28679
rect 27580 28648 28825 28676
rect 27580 28636 27586 28648
rect 28813 28645 28825 28648
rect 28859 28676 28871 28679
rect 29914 28676 29920 28688
rect 28859 28648 29920 28676
rect 28859 28645 28871 28648
rect 28813 28639 28871 28645
rect 29914 28636 29920 28648
rect 29972 28636 29978 28688
rect 30006 28636 30012 28688
rect 30064 28676 30070 28688
rect 30742 28676 30748 28688
rect 30064 28648 30748 28676
rect 30064 28636 30070 28648
rect 30742 28636 30748 28648
rect 30800 28636 30806 28688
rect 29730 28608 29736 28620
rect 24596 28580 29736 28608
rect 23293 28571 23351 28577
rect 29730 28568 29736 28580
rect 29788 28568 29794 28620
rect 22051 28543 22109 28549
rect 22051 28540 22063 28543
rect 21600 28512 22063 28540
rect 21600 28500 21606 28512
rect 22051 28509 22063 28512
rect 22097 28509 22109 28543
rect 22051 28503 22109 28509
rect 22189 28543 22247 28549
rect 22189 28509 22201 28543
rect 22235 28509 22247 28543
rect 22189 28503 22247 28509
rect 22281 28543 22339 28549
rect 22281 28509 22293 28543
rect 22327 28509 22339 28543
rect 22281 28503 22339 28509
rect 22462 28500 22468 28552
rect 22520 28540 22526 28552
rect 25317 28543 25375 28549
rect 25317 28540 25329 28543
rect 22520 28512 22613 28540
rect 22940 28512 25329 28540
rect 22520 28500 22526 28512
rect 22480 28472 22508 28500
rect 22940 28484 22968 28512
rect 25317 28509 25329 28512
rect 25363 28540 25375 28543
rect 27801 28543 27859 28549
rect 25363 28512 27743 28540
rect 25363 28509 25375 28512
rect 25317 28503 25375 28509
rect 22922 28472 22928 28484
rect 21376 28444 22508 28472
rect 22883 28444 22928 28472
rect 22922 28432 22928 28444
rect 22980 28432 22986 28484
rect 23109 28475 23167 28481
rect 23109 28441 23121 28475
rect 23155 28441 23167 28475
rect 23109 28435 23167 28441
rect 17129 28407 17187 28413
rect 17129 28404 17141 28407
rect 16816 28376 17141 28404
rect 16816 28364 16822 28376
rect 17129 28373 17141 28376
rect 17175 28373 17187 28407
rect 18248 28404 18276 28432
rect 18598 28404 18604 28416
rect 18248 28376 18604 28404
rect 17129 28367 17187 28373
rect 18598 28364 18604 28376
rect 18656 28364 18662 28416
rect 19058 28364 19064 28416
rect 19116 28404 19122 28416
rect 19426 28404 19432 28416
rect 19116 28376 19432 28404
rect 19116 28364 19122 28376
rect 19426 28364 19432 28376
rect 19484 28364 19490 28416
rect 20990 28364 20996 28416
rect 21048 28404 21054 28416
rect 21174 28404 21180 28416
rect 21048 28376 21180 28404
rect 21048 28364 21054 28376
rect 21174 28364 21180 28376
rect 21232 28364 21238 28416
rect 21818 28364 21824 28416
rect 21876 28404 21882 28416
rect 23124 28404 23152 28435
rect 23290 28432 23296 28484
rect 23348 28472 23354 28484
rect 24397 28475 24455 28481
rect 24397 28472 24409 28475
rect 23348 28444 24409 28472
rect 23348 28432 23354 28444
rect 24397 28441 24409 28444
rect 24443 28441 24455 28475
rect 24397 28435 24455 28441
rect 25501 28475 25559 28481
rect 25501 28441 25513 28475
rect 25547 28472 25559 28475
rect 25590 28472 25596 28484
rect 25547 28444 25596 28472
rect 25547 28441 25559 28444
rect 25501 28435 25559 28441
rect 25590 28432 25596 28444
rect 25648 28432 25654 28484
rect 26970 28472 26976 28484
rect 26931 28444 26976 28472
rect 26970 28432 26976 28444
rect 27028 28432 27034 28484
rect 27715 28472 27743 28512
rect 27801 28509 27813 28543
rect 27847 28540 27859 28543
rect 27890 28540 27896 28552
rect 27847 28512 27896 28540
rect 27847 28509 27859 28512
rect 27801 28503 27859 28509
rect 27890 28500 27896 28512
rect 27948 28500 27954 28552
rect 28074 28540 28080 28552
rect 28035 28512 28080 28540
rect 28074 28500 28080 28512
rect 28132 28500 28138 28552
rect 30006 28540 30012 28552
rect 29967 28512 30012 28540
rect 30006 28500 30012 28512
rect 30064 28500 30070 28552
rect 30101 28543 30159 28549
rect 30101 28509 30113 28543
rect 30147 28509 30159 28543
rect 30101 28503 30159 28509
rect 27715 28444 28120 28472
rect 21876 28376 23152 28404
rect 21876 28364 21882 28376
rect 23474 28364 23480 28416
rect 23532 28404 23538 28416
rect 24210 28404 24216 28416
rect 23532 28376 24216 28404
rect 23532 28364 23538 28376
rect 24210 28364 24216 28376
rect 24268 28364 24274 28416
rect 24486 28364 24492 28416
rect 24544 28404 24550 28416
rect 24597 28407 24655 28413
rect 24597 28404 24609 28407
rect 24544 28376 24609 28404
rect 24544 28364 24550 28376
rect 24597 28373 24609 28376
rect 24643 28373 24655 28407
rect 24762 28404 24768 28416
rect 24723 28376 24768 28404
rect 24597 28367 24655 28373
rect 24762 28364 24768 28376
rect 24820 28364 24826 28416
rect 26786 28364 26792 28416
rect 26844 28404 26850 28416
rect 27065 28407 27123 28413
rect 27065 28404 27077 28407
rect 26844 28376 27077 28404
rect 26844 28364 26850 28376
rect 27065 28373 27077 28376
rect 27111 28373 27123 28407
rect 27982 28404 27988 28416
rect 27943 28376 27988 28404
rect 27065 28367 27123 28373
rect 27982 28364 27988 28376
rect 28040 28364 28046 28416
rect 28092 28404 28120 28444
rect 28350 28432 28356 28484
rect 28408 28472 28414 28484
rect 28629 28475 28687 28481
rect 28629 28472 28641 28475
rect 28408 28444 28641 28472
rect 28408 28432 28414 28444
rect 28629 28441 28641 28444
rect 28675 28441 28687 28475
rect 28629 28435 28687 28441
rect 29822 28432 29828 28484
rect 29880 28472 29886 28484
rect 30116 28472 30144 28503
rect 30190 28500 30196 28552
rect 30248 28540 30254 28552
rect 30377 28543 30435 28549
rect 30248 28512 30293 28540
rect 30248 28500 30254 28512
rect 30377 28509 30389 28543
rect 30423 28509 30435 28543
rect 30377 28503 30435 28509
rect 29880 28444 30144 28472
rect 29880 28432 29886 28444
rect 28994 28404 29000 28416
rect 28092 28376 29000 28404
rect 28994 28364 29000 28376
rect 29052 28364 29058 28416
rect 29914 28364 29920 28416
rect 29972 28404 29978 28416
rect 30392 28404 30420 28503
rect 31110 28472 31116 28484
rect 31071 28444 31116 28472
rect 31110 28432 31116 28444
rect 31168 28432 31174 28484
rect 29972 28376 30420 28404
rect 29972 28364 29978 28376
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 6362 28160 6368 28212
rect 6420 28200 6426 28212
rect 6641 28203 6699 28209
rect 6641 28200 6653 28203
rect 6420 28172 6653 28200
rect 6420 28160 6426 28172
rect 6641 28169 6653 28172
rect 6687 28169 6699 28203
rect 8662 28200 8668 28212
rect 8623 28172 8668 28200
rect 6641 28163 6699 28169
rect 8662 28160 8668 28172
rect 8720 28160 8726 28212
rect 10778 28160 10784 28212
rect 10836 28200 10842 28212
rect 10836 28172 12434 28200
rect 10836 28160 10842 28172
rect 12406 28132 12434 28172
rect 13538 28160 13544 28212
rect 13596 28200 13602 28212
rect 13633 28203 13691 28209
rect 13633 28200 13645 28203
rect 13596 28172 13645 28200
rect 13596 28160 13602 28172
rect 13633 28169 13645 28172
rect 13679 28169 13691 28203
rect 15470 28200 15476 28212
rect 15431 28172 15476 28200
rect 13633 28163 13691 28169
rect 15470 28160 15476 28172
rect 15528 28160 15534 28212
rect 18046 28160 18052 28212
rect 18104 28200 18110 28212
rect 18233 28203 18291 28209
rect 18233 28200 18245 28203
rect 18104 28172 18245 28200
rect 18104 28160 18110 28172
rect 18233 28169 18245 28172
rect 18279 28169 18291 28203
rect 19058 28200 19064 28212
rect 19019 28172 19064 28200
rect 18233 28163 18291 28169
rect 19058 28160 19064 28172
rect 19116 28160 19122 28212
rect 20898 28160 20904 28212
rect 20956 28200 20962 28212
rect 21177 28203 21235 28209
rect 21177 28200 21189 28203
rect 20956 28172 21189 28200
rect 20956 28160 20962 28172
rect 21177 28169 21189 28172
rect 21223 28169 21235 28203
rect 21177 28163 21235 28169
rect 26326 28160 26332 28212
rect 26384 28200 26390 28212
rect 26421 28203 26479 28209
rect 26421 28200 26433 28203
rect 26384 28172 26433 28200
rect 26384 28160 26390 28172
rect 26421 28169 26433 28172
rect 26467 28169 26479 28203
rect 26421 28163 26479 28169
rect 28994 28160 29000 28212
rect 29052 28200 29058 28212
rect 31018 28200 31024 28212
rect 29052 28172 30696 28200
rect 30979 28172 31024 28200
rect 29052 28160 29058 28172
rect 16758 28132 16764 28144
rect 7300 28104 9076 28132
rect 12406 28104 13584 28132
rect 6825 28067 6883 28073
rect 6825 28033 6837 28067
rect 6871 28064 6883 28067
rect 7190 28064 7196 28076
rect 6871 28036 7196 28064
rect 6871 28033 6883 28036
rect 6825 28027 6883 28033
rect 7190 28024 7196 28036
rect 7248 28024 7254 28076
rect 7300 28073 7328 28104
rect 9048 28076 9076 28104
rect 7558 28073 7564 28076
rect 7285 28067 7343 28073
rect 7285 28033 7297 28067
rect 7331 28033 7343 28067
rect 7552 28064 7564 28073
rect 7519 28036 7564 28064
rect 7285 28027 7343 28033
rect 7552 28027 7564 28036
rect 7558 28024 7564 28027
rect 7616 28024 7622 28076
rect 9030 28024 9036 28076
rect 9088 28064 9094 28076
rect 9125 28067 9183 28073
rect 9125 28064 9137 28067
rect 9088 28036 9137 28064
rect 9088 28024 9094 28036
rect 9125 28033 9137 28036
rect 9171 28033 9183 28067
rect 9125 28027 9183 28033
rect 9214 28024 9220 28076
rect 9272 28064 9278 28076
rect 9381 28067 9439 28073
rect 9381 28064 9393 28067
rect 9272 28036 9393 28064
rect 9272 28024 9278 28036
rect 9381 28033 9393 28036
rect 9427 28033 9439 28067
rect 11514 28064 11520 28076
rect 11475 28036 11520 28064
rect 9381 28027 9439 28033
rect 11514 28024 11520 28036
rect 11572 28024 11578 28076
rect 11606 28024 11612 28076
rect 11664 28064 11670 28076
rect 13556 28073 13584 28104
rect 15764 28104 16764 28132
rect 11773 28067 11831 28073
rect 11773 28064 11785 28067
rect 11664 28036 11785 28064
rect 11664 28024 11670 28036
rect 11773 28033 11785 28036
rect 11819 28033 11831 28067
rect 11773 28027 11831 28033
rect 13541 28067 13599 28073
rect 13541 28033 13553 28067
rect 13587 28064 13599 28067
rect 14829 28067 14887 28073
rect 14829 28064 14841 28067
rect 13587 28036 14841 28064
rect 13587 28033 13599 28036
rect 13541 28027 13599 28033
rect 14829 28033 14841 28036
rect 14875 28064 14887 28067
rect 14918 28064 14924 28076
rect 14875 28036 14924 28064
rect 14875 28033 14887 28036
rect 14829 28027 14887 28033
rect 14918 28024 14924 28036
rect 14976 28024 14982 28076
rect 15764 28073 15792 28104
rect 16758 28092 16764 28104
rect 16816 28092 16822 28144
rect 19426 28132 19432 28144
rect 16868 28104 17632 28132
rect 15749 28067 15807 28073
rect 15749 28033 15761 28067
rect 15795 28033 15807 28067
rect 15749 28027 15807 28033
rect 15841 28067 15899 28073
rect 15841 28033 15853 28067
rect 15887 28033 15899 28067
rect 15841 28027 15899 28033
rect 15954 28067 16012 28073
rect 15954 28033 15966 28067
rect 16000 28064 16012 28067
rect 16000 28036 16068 28064
rect 16000 28033 16012 28036
rect 15954 28027 16012 28033
rect 15010 27956 15016 28008
rect 15068 27996 15074 28008
rect 15856 27996 15884 28027
rect 15068 27968 15884 27996
rect 16040 27996 16068 28036
rect 16114 28024 16120 28076
rect 16172 28064 16178 28076
rect 16868 28073 16896 28104
rect 16853 28067 16911 28073
rect 16172 28036 16217 28064
rect 16172 28024 16178 28036
rect 16853 28033 16865 28067
rect 16899 28033 16911 28067
rect 16853 28027 16911 28033
rect 17120 28067 17178 28073
rect 17120 28033 17132 28067
rect 17166 28064 17178 28067
rect 17494 28064 17500 28076
rect 17166 28036 17500 28064
rect 17166 28033 17178 28036
rect 17120 28027 17178 28033
rect 17494 28024 17500 28036
rect 17552 28024 17558 28076
rect 17604 28064 17632 28104
rect 18540 28104 19432 28132
rect 18540 28064 18568 28104
rect 19426 28092 19432 28104
rect 19484 28092 19490 28144
rect 19889 28135 19947 28141
rect 19889 28101 19901 28135
rect 19935 28132 19947 28135
rect 19978 28132 19984 28144
rect 19935 28104 19984 28132
rect 19935 28101 19947 28104
rect 19889 28095 19947 28101
rect 19978 28092 19984 28104
rect 20036 28092 20042 28144
rect 24210 28132 24216 28144
rect 24171 28104 24216 28132
rect 24210 28092 24216 28104
rect 24268 28092 24274 28144
rect 27341 28135 27399 28141
rect 27341 28101 27353 28135
rect 27387 28132 27399 28135
rect 30374 28132 30380 28144
rect 27387 28104 30380 28132
rect 27387 28101 27399 28104
rect 27341 28095 27399 28101
rect 30374 28092 30380 28104
rect 30432 28132 30438 28144
rect 30432 28104 30604 28132
rect 30432 28092 30438 28104
rect 17604 28036 18568 28064
rect 18598 28024 18604 28076
rect 18656 28064 18662 28076
rect 18877 28067 18935 28073
rect 18877 28064 18889 28067
rect 18656 28036 18889 28064
rect 18656 28024 18662 28036
rect 18877 28033 18889 28036
rect 18923 28033 18935 28067
rect 18877 28027 18935 28033
rect 19705 28067 19763 28073
rect 19705 28033 19717 28067
rect 19751 28064 19763 28067
rect 20254 28064 20260 28076
rect 19751 28036 20260 28064
rect 19751 28033 19763 28036
rect 19705 28027 19763 28033
rect 16298 27996 16304 28008
rect 16040 27968 16304 27996
rect 15068 27956 15074 27968
rect 16298 27956 16304 27968
rect 16356 27956 16362 28008
rect 17862 27956 17868 28008
rect 17920 27996 17926 28008
rect 19720 27996 19748 28027
rect 20254 28024 20260 28036
rect 20312 28024 20318 28076
rect 20990 28064 20996 28076
rect 20951 28036 20996 28064
rect 20990 28024 20996 28036
rect 21048 28024 21054 28076
rect 21910 28064 21916 28076
rect 21871 28036 21916 28064
rect 21910 28024 21916 28036
rect 21968 28024 21974 28076
rect 22186 28073 22192 28076
rect 22180 28027 22192 28073
rect 22244 28064 22250 28076
rect 25038 28064 25044 28076
rect 22244 28036 22280 28064
rect 24999 28036 25044 28064
rect 22186 28024 22192 28027
rect 22244 28024 22250 28036
rect 25038 28024 25044 28036
rect 25096 28024 25102 28076
rect 25314 28073 25320 28076
rect 25308 28027 25320 28073
rect 25372 28064 25378 28076
rect 25372 28036 25408 28064
rect 25314 28024 25320 28027
rect 25372 28024 25378 28036
rect 26970 28024 26976 28076
rect 27028 28064 27034 28076
rect 28350 28064 28356 28076
rect 27028 28036 28356 28064
rect 27028 28024 27034 28036
rect 28350 28024 28356 28036
rect 28408 28024 28414 28076
rect 29638 28024 29644 28076
rect 29696 28064 29702 28076
rect 29779 28067 29837 28073
rect 29779 28064 29791 28067
rect 29696 28036 29791 28064
rect 29696 28024 29702 28036
rect 29779 28033 29791 28036
rect 29825 28033 29837 28067
rect 29914 28064 29920 28076
rect 29875 28036 29920 28064
rect 29779 28027 29837 28033
rect 29914 28024 29920 28036
rect 29972 28024 29978 28076
rect 30009 28070 30067 28076
rect 30009 28036 30021 28070
rect 30055 28036 30067 28070
rect 30190 28064 30196 28076
rect 30151 28036 30196 28064
rect 30009 28030 30067 28036
rect 17920 27968 19748 27996
rect 20809 27999 20867 28005
rect 17920 27956 17926 27968
rect 20809 27965 20821 27999
rect 20855 27996 20867 27999
rect 21542 27996 21548 28008
rect 20855 27968 21548 27996
rect 20855 27965 20867 27968
rect 20809 27959 20867 27965
rect 21542 27956 21548 27968
rect 21600 27956 21606 28008
rect 28994 27956 29000 28008
rect 29052 27996 29058 28008
rect 30024 27996 30052 28030
rect 30190 28024 30196 28036
rect 30248 28024 30254 28076
rect 29052 27968 30052 27996
rect 30576 27996 30604 28104
rect 30668 28073 30696 28172
rect 31018 28160 31024 28172
rect 31076 28160 31082 28212
rect 31110 28132 31116 28144
rect 30760 28104 31116 28132
rect 30653 28067 30711 28073
rect 30653 28033 30665 28067
rect 30699 28033 30711 28067
rect 30653 28027 30711 28033
rect 30760 27996 30788 28104
rect 31110 28092 31116 28104
rect 31168 28092 31174 28144
rect 30837 28067 30895 28073
rect 30837 28033 30849 28067
rect 30883 28033 30895 28067
rect 30837 28027 30895 28033
rect 30576 27968 30788 27996
rect 29052 27956 29058 27968
rect 12710 27888 12716 27940
rect 12768 27928 12774 27940
rect 12897 27931 12955 27937
rect 12897 27928 12909 27931
rect 12768 27900 12909 27928
rect 12768 27888 12774 27900
rect 12897 27897 12909 27900
rect 12943 27928 12955 27931
rect 16666 27928 16672 27940
rect 12943 27900 16672 27928
rect 12943 27897 12955 27900
rect 12897 27891 12955 27897
rect 16666 27888 16672 27900
rect 16724 27888 16730 27940
rect 19242 27888 19248 27940
rect 19300 27928 19306 27940
rect 19886 27928 19892 27940
rect 19300 27900 19892 27928
rect 19300 27888 19306 27900
rect 19886 27888 19892 27900
rect 19944 27888 19950 27940
rect 23293 27931 23351 27937
rect 23293 27897 23305 27931
rect 23339 27928 23351 27931
rect 23382 27928 23388 27940
rect 23339 27900 23388 27928
rect 23339 27897 23351 27900
rect 23293 27891 23351 27897
rect 10502 27860 10508 27872
rect 10463 27832 10508 27860
rect 10502 27820 10508 27832
rect 10560 27820 10566 27872
rect 14366 27820 14372 27872
rect 14424 27860 14430 27872
rect 14921 27863 14979 27869
rect 14921 27860 14933 27863
rect 14424 27832 14933 27860
rect 14424 27820 14430 27832
rect 14921 27829 14933 27832
rect 14967 27860 14979 27863
rect 19260 27860 19288 27888
rect 14967 27832 19288 27860
rect 14967 27829 14979 27832
rect 14921 27823 14979 27829
rect 19334 27820 19340 27872
rect 19392 27860 19398 27872
rect 19518 27860 19524 27872
rect 19392 27832 19524 27860
rect 19392 27820 19398 27832
rect 19518 27820 19524 27832
rect 19576 27860 19582 27872
rect 20162 27860 20168 27872
rect 19576 27832 20168 27860
rect 19576 27820 19582 27832
rect 20162 27820 20168 27832
rect 20220 27820 20226 27872
rect 20438 27820 20444 27872
rect 20496 27860 20502 27872
rect 20622 27860 20628 27872
rect 20496 27832 20628 27860
rect 20496 27820 20502 27832
rect 20622 27820 20628 27832
rect 20680 27820 20686 27872
rect 20898 27820 20904 27872
rect 20956 27860 20962 27872
rect 23308 27860 23336 27891
rect 23382 27888 23388 27900
rect 23440 27888 23446 27940
rect 23842 27928 23848 27940
rect 23803 27900 23848 27928
rect 23842 27888 23848 27900
rect 23900 27888 23906 27940
rect 24762 27928 24768 27940
rect 24228 27900 24768 27928
rect 24228 27869 24256 27900
rect 24762 27888 24768 27900
rect 24820 27888 24826 27940
rect 29454 27888 29460 27940
rect 29512 27928 29518 27940
rect 30852 27928 30880 28027
rect 29512 27900 30880 27928
rect 29512 27888 29518 27900
rect 20956 27832 23336 27860
rect 24213 27863 24271 27869
rect 20956 27820 20962 27832
rect 24213 27829 24225 27863
rect 24259 27829 24271 27863
rect 24213 27823 24271 27829
rect 24302 27820 24308 27872
rect 24360 27860 24366 27872
rect 24397 27863 24455 27869
rect 24397 27860 24409 27863
rect 24360 27832 24409 27860
rect 24360 27820 24366 27832
rect 24397 27829 24409 27832
rect 24443 27829 24455 27863
rect 24397 27823 24455 27829
rect 27614 27820 27620 27872
rect 27672 27860 27678 27872
rect 28629 27863 28687 27869
rect 28629 27860 28641 27863
rect 27672 27832 28641 27860
rect 27672 27820 27678 27832
rect 28629 27829 28641 27832
rect 28675 27829 28687 27863
rect 28629 27823 28687 27829
rect 29549 27863 29607 27869
rect 29549 27829 29561 27863
rect 29595 27860 29607 27863
rect 30282 27860 30288 27872
rect 29595 27832 30288 27860
rect 29595 27829 29607 27832
rect 29549 27823 29607 27829
rect 30282 27820 30288 27832
rect 30340 27820 30346 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 6546 27616 6552 27668
rect 6604 27656 6610 27668
rect 6733 27659 6791 27665
rect 6733 27656 6745 27659
rect 6604 27628 6745 27656
rect 6604 27616 6610 27628
rect 6733 27625 6745 27628
rect 6779 27625 6791 27659
rect 6733 27619 6791 27625
rect 7929 27659 7987 27665
rect 7929 27625 7941 27659
rect 7975 27656 7987 27659
rect 10502 27656 10508 27668
rect 7975 27628 10508 27656
rect 7975 27625 7987 27628
rect 7929 27619 7987 27625
rect 10502 27616 10508 27628
rect 10560 27616 10566 27668
rect 11241 27659 11299 27665
rect 11241 27625 11253 27659
rect 11287 27656 11299 27659
rect 11606 27656 11612 27668
rect 11287 27628 11612 27656
rect 11287 27625 11299 27628
rect 11241 27619 11299 27625
rect 11606 27616 11612 27628
rect 11664 27616 11670 27668
rect 17494 27656 17500 27668
rect 15396 27628 16344 27656
rect 17455 27628 17500 27656
rect 10689 27591 10747 27597
rect 10689 27557 10701 27591
rect 10735 27588 10747 27591
rect 10870 27588 10876 27600
rect 10735 27560 10876 27588
rect 10735 27557 10747 27560
rect 10689 27551 10747 27557
rect 10870 27548 10876 27560
rect 10928 27548 10934 27600
rect 14274 27588 14280 27600
rect 11624 27560 14280 27588
rect 5353 27455 5411 27461
rect 5353 27421 5365 27455
rect 5399 27452 5411 27455
rect 5442 27452 5448 27464
rect 5399 27424 5448 27452
rect 5399 27421 5411 27424
rect 5353 27415 5411 27421
rect 5442 27412 5448 27424
rect 5500 27412 5506 27464
rect 5620 27455 5678 27461
rect 5620 27421 5632 27455
rect 5666 27452 5678 27455
rect 5902 27452 5908 27464
rect 5666 27424 5908 27452
rect 5666 27421 5678 27424
rect 5620 27415 5678 27421
rect 5902 27412 5908 27424
rect 5960 27412 5966 27464
rect 9950 27412 9956 27464
rect 10008 27452 10014 27464
rect 10505 27455 10563 27461
rect 10505 27452 10517 27455
rect 10008 27424 10517 27452
rect 10008 27412 10014 27424
rect 10505 27421 10517 27424
rect 10551 27452 10563 27455
rect 10778 27452 10784 27464
rect 10551 27424 10784 27452
rect 10551 27421 10563 27424
rect 10505 27415 10563 27421
rect 10778 27412 10784 27424
rect 10836 27412 10842 27464
rect 11422 27412 11428 27464
rect 11480 27452 11486 27464
rect 11624 27461 11652 27560
rect 14274 27548 14280 27560
rect 14332 27548 14338 27600
rect 15396 27588 15424 27628
rect 14568 27560 15424 27588
rect 16316 27588 16344 27628
rect 17494 27616 17500 27628
rect 17552 27616 17558 27668
rect 19058 27656 19064 27668
rect 17604 27628 19064 27656
rect 16758 27588 16764 27600
rect 16316 27560 16436 27588
rect 16671 27560 16764 27588
rect 12805 27523 12863 27529
rect 12805 27520 12817 27523
rect 11716 27492 12817 27520
rect 11716 27461 11744 27492
rect 12805 27489 12817 27492
rect 12851 27489 12863 27523
rect 14568 27520 14596 27560
rect 12805 27483 12863 27489
rect 13280 27492 14596 27520
rect 11517 27455 11575 27461
rect 11517 27452 11529 27455
rect 11480 27424 11529 27452
rect 11480 27412 11486 27424
rect 11517 27421 11529 27424
rect 11563 27421 11575 27455
rect 11517 27415 11575 27421
rect 11609 27455 11667 27461
rect 11609 27421 11621 27455
rect 11655 27421 11667 27455
rect 11609 27415 11667 27421
rect 11701 27455 11759 27461
rect 11701 27421 11713 27455
rect 11747 27421 11759 27455
rect 11882 27452 11888 27464
rect 11843 27424 11888 27452
rect 11701 27415 11759 27421
rect 7742 27384 7748 27396
rect 7703 27356 7748 27384
rect 7742 27344 7748 27356
rect 7800 27344 7806 27396
rect 7926 27344 7932 27396
rect 7984 27393 7990 27396
rect 7984 27387 8003 27393
rect 7991 27353 8003 27387
rect 7984 27347 8003 27353
rect 7984 27344 7990 27347
rect 9858 27344 9864 27396
rect 9916 27384 9922 27396
rect 11624 27384 11652 27415
rect 11882 27412 11888 27424
rect 11940 27412 11946 27464
rect 12621 27455 12679 27461
rect 12621 27421 12633 27455
rect 12667 27452 12679 27455
rect 12710 27452 12716 27464
rect 12667 27424 12716 27452
rect 12667 27421 12679 27424
rect 12621 27415 12679 27421
rect 12710 27412 12716 27424
rect 12768 27412 12774 27464
rect 13280 27461 13308 27492
rect 14642 27480 14648 27532
rect 14700 27520 14706 27532
rect 16408 27520 16436 27560
rect 16758 27548 16764 27560
rect 16816 27588 16822 27600
rect 17402 27588 17408 27600
rect 16816 27560 17408 27588
rect 16816 27548 16822 27560
rect 17402 27548 17408 27560
rect 17460 27548 17466 27600
rect 17604 27520 17632 27628
rect 19058 27616 19064 27628
rect 19116 27616 19122 27668
rect 19886 27656 19892 27668
rect 19720 27628 19892 27656
rect 19720 27600 19748 27628
rect 19886 27616 19892 27628
rect 19944 27616 19950 27668
rect 20990 27616 20996 27668
rect 21048 27656 21054 27668
rect 24026 27656 24032 27668
rect 21048 27628 24032 27656
rect 21048 27616 21054 27628
rect 24026 27616 24032 27628
rect 24084 27616 24090 27668
rect 26786 27616 26792 27668
rect 26844 27656 26850 27668
rect 30190 27656 30196 27668
rect 26844 27628 30196 27656
rect 26844 27616 26850 27628
rect 30190 27616 30196 27628
rect 30248 27616 30254 27668
rect 19334 27588 19340 27600
rect 14700 27492 15516 27520
rect 16408 27492 17632 27520
rect 17696 27560 19340 27588
rect 14700 27480 14706 27492
rect 13265 27455 13323 27461
rect 13265 27421 13277 27455
rect 13311 27421 13323 27455
rect 13265 27415 13323 27421
rect 9916 27356 11652 27384
rect 12437 27387 12495 27393
rect 9916 27344 9922 27356
rect 12437 27353 12449 27387
rect 12483 27384 12495 27387
rect 13170 27384 13176 27396
rect 12483 27356 13176 27384
rect 12483 27353 12495 27356
rect 12437 27347 12495 27353
rect 13170 27344 13176 27356
rect 13228 27344 13234 27396
rect 8110 27316 8116 27328
rect 8071 27288 8116 27316
rect 8110 27276 8116 27288
rect 8168 27276 8174 27328
rect 9306 27276 9312 27328
rect 9364 27316 9370 27328
rect 13280 27316 13308 27415
rect 14090 27412 14096 27464
rect 14148 27452 14154 27464
rect 15381 27455 15439 27461
rect 15381 27452 15393 27455
rect 14148 27424 15393 27452
rect 14148 27412 14154 27424
rect 15381 27421 15393 27424
rect 15427 27421 15439 27455
rect 15488 27452 15516 27492
rect 17696 27461 17724 27560
rect 19334 27548 19340 27560
rect 19392 27548 19398 27600
rect 19702 27548 19708 27600
rect 19760 27548 19766 27600
rect 21545 27591 21603 27597
rect 21545 27557 21557 27591
rect 21591 27588 21603 27591
rect 22186 27588 22192 27600
rect 21591 27560 22192 27588
rect 21591 27557 21603 27560
rect 21545 27551 21603 27557
rect 22186 27548 22192 27560
rect 22244 27548 22250 27600
rect 23290 27588 23296 27600
rect 22848 27560 23296 27588
rect 21085 27523 21143 27529
rect 17926 27492 19656 27520
rect 17681 27455 17739 27461
rect 15488 27424 17632 27452
rect 15381 27415 15439 27421
rect 14366 27344 14372 27396
rect 14424 27384 14430 27396
rect 14553 27387 14611 27393
rect 14553 27384 14565 27387
rect 14424 27356 14565 27384
rect 14424 27344 14430 27356
rect 14553 27353 14565 27356
rect 14599 27353 14611 27387
rect 14553 27347 14611 27353
rect 14737 27387 14795 27393
rect 14737 27353 14749 27387
rect 14783 27384 14795 27387
rect 14826 27384 14832 27396
rect 14783 27356 14832 27384
rect 14783 27353 14795 27356
rect 14737 27347 14795 27353
rect 14826 27344 14832 27356
rect 14884 27384 14890 27396
rect 15286 27384 15292 27396
rect 14884 27356 15292 27384
rect 14884 27344 14890 27356
rect 15286 27344 15292 27356
rect 15344 27344 15350 27396
rect 15470 27344 15476 27396
rect 15528 27384 15534 27396
rect 15626 27387 15684 27393
rect 15626 27384 15638 27387
rect 15528 27356 15638 27384
rect 15528 27344 15534 27356
rect 15626 27353 15638 27356
rect 15672 27353 15684 27387
rect 17604 27384 17632 27424
rect 17681 27421 17693 27455
rect 17727 27421 17739 27455
rect 17681 27415 17739 27421
rect 17926 27384 17954 27492
rect 19518 27452 19524 27464
rect 19479 27424 19524 27452
rect 19518 27412 19524 27424
rect 19576 27412 19582 27464
rect 19628 27461 19656 27492
rect 20640 27492 21036 27520
rect 19613 27455 19671 27461
rect 19613 27421 19625 27455
rect 19659 27421 19671 27455
rect 19613 27415 19671 27421
rect 17604 27356 17954 27384
rect 15626 27347 15684 27353
rect 18966 27344 18972 27396
rect 19024 27384 19030 27396
rect 19625 27384 19653 27415
rect 19702 27412 19708 27464
rect 19760 27452 19766 27464
rect 19889 27455 19947 27461
rect 19760 27424 19805 27452
rect 19760 27412 19766 27424
rect 19889 27421 19901 27455
rect 19935 27452 19947 27455
rect 20254 27452 20260 27464
rect 19935 27424 20260 27452
rect 19935 27421 19947 27424
rect 19889 27415 19947 27421
rect 20254 27412 20260 27424
rect 20312 27412 20318 27464
rect 20640 27384 20668 27492
rect 20898 27452 20904 27464
rect 20859 27424 20904 27452
rect 20898 27412 20904 27424
rect 20956 27412 20962 27464
rect 21008 27452 21036 27492
rect 21085 27489 21097 27523
rect 21131 27520 21143 27523
rect 21131 27492 22048 27520
rect 21131 27489 21143 27492
rect 21085 27483 21143 27489
rect 21266 27452 21272 27464
rect 21008 27424 21272 27452
rect 21266 27412 21272 27424
rect 21324 27412 21330 27464
rect 21358 27412 21364 27464
rect 21416 27452 21422 27464
rect 21818 27452 21824 27464
rect 21416 27424 21824 27452
rect 21416 27412 21422 27424
rect 21818 27412 21824 27424
rect 21876 27412 21882 27464
rect 22020 27461 22048 27492
rect 21913 27455 21971 27461
rect 21913 27421 21925 27455
rect 21959 27421 21971 27455
rect 21913 27415 21971 27421
rect 22005 27455 22063 27461
rect 22005 27421 22017 27455
rect 22051 27421 22063 27455
rect 22005 27415 22063 27421
rect 22189 27455 22247 27461
rect 22189 27421 22201 27455
rect 22235 27421 22247 27455
rect 22189 27415 22247 27421
rect 19024 27356 19380 27384
rect 19625 27356 20668 27384
rect 20717 27387 20775 27393
rect 19024 27344 19030 27356
rect 9364 27288 13308 27316
rect 13449 27319 13507 27325
rect 9364 27276 9370 27288
rect 13449 27285 13461 27319
rect 13495 27316 13507 27319
rect 13538 27316 13544 27328
rect 13495 27288 13544 27316
rect 13495 27285 13507 27288
rect 13449 27279 13507 27285
rect 13538 27276 13544 27288
rect 13596 27316 13602 27328
rect 13814 27316 13820 27328
rect 13596 27288 13820 27316
rect 13596 27276 13602 27288
rect 13814 27276 13820 27288
rect 13872 27276 13878 27328
rect 14921 27319 14979 27325
rect 14921 27285 14933 27319
rect 14967 27316 14979 27319
rect 15838 27316 15844 27328
rect 14967 27288 15844 27316
rect 14967 27285 14979 27288
rect 14921 27279 14979 27285
rect 15838 27276 15844 27288
rect 15896 27276 15902 27328
rect 19242 27316 19248 27328
rect 19203 27288 19248 27316
rect 19242 27276 19248 27288
rect 19300 27276 19306 27328
rect 19352 27316 19380 27356
rect 20717 27353 20729 27387
rect 20763 27353 20775 27387
rect 21284 27384 21312 27412
rect 21928 27384 21956 27415
rect 21284 27356 21956 27384
rect 22204 27384 22232 27415
rect 22278 27412 22284 27464
rect 22336 27452 22342 27464
rect 22848 27461 22876 27560
rect 23290 27548 23296 27560
rect 23348 27548 23354 27600
rect 23842 27548 23848 27600
rect 23900 27588 23906 27600
rect 24673 27591 24731 27597
rect 24673 27588 24685 27591
rect 23900 27560 24685 27588
rect 23900 27548 23906 27560
rect 24673 27557 24685 27560
rect 24719 27557 24731 27591
rect 24673 27551 24731 27557
rect 26421 27591 26479 27597
rect 26421 27557 26433 27591
rect 26467 27588 26479 27591
rect 27522 27588 27528 27600
rect 26467 27560 27528 27588
rect 26467 27557 26479 27560
rect 26421 27551 26479 27557
rect 27522 27548 27528 27560
rect 27580 27548 27586 27600
rect 27890 27548 27896 27600
rect 27948 27588 27954 27600
rect 28258 27588 28264 27600
rect 27948 27560 28264 27588
rect 27948 27548 27954 27560
rect 28258 27548 28264 27560
rect 28316 27588 28322 27600
rect 28316 27560 29408 27588
rect 28316 27548 28322 27560
rect 23198 27480 23204 27532
rect 23256 27520 23262 27532
rect 28534 27520 28540 27532
rect 23256 27492 24256 27520
rect 23256 27480 23262 27492
rect 22833 27455 22891 27461
rect 22833 27452 22845 27455
rect 22336 27424 22845 27452
rect 22336 27412 22342 27424
rect 22833 27421 22845 27424
rect 22879 27421 22891 27455
rect 22833 27415 22891 27421
rect 23014 27412 23020 27464
rect 23072 27452 23078 27464
rect 24228 27452 24256 27492
rect 25792 27492 27614 27520
rect 25792 27461 25820 27492
rect 25777 27455 25835 27461
rect 23072 27424 24164 27452
rect 24228 27424 24532 27452
rect 23072 27412 23078 27424
rect 23290 27384 23296 27396
rect 22204 27356 23296 27384
rect 20717 27347 20775 27353
rect 20732 27316 20760 27347
rect 23290 27344 23296 27356
rect 23348 27344 23354 27396
rect 23661 27387 23719 27393
rect 23661 27353 23673 27387
rect 23707 27384 23719 27387
rect 24026 27384 24032 27396
rect 23707 27356 24032 27384
rect 23707 27353 23719 27356
rect 23661 27347 23719 27353
rect 24026 27344 24032 27356
rect 24084 27344 24090 27396
rect 22278 27316 22284 27328
rect 19352 27288 22284 27316
rect 22278 27276 22284 27288
rect 22336 27276 22342 27328
rect 23017 27319 23075 27325
rect 23017 27285 23029 27319
rect 23063 27316 23075 27319
rect 23474 27316 23480 27328
rect 23063 27288 23480 27316
rect 23063 27285 23075 27288
rect 23017 27279 23075 27285
rect 23474 27276 23480 27288
rect 23532 27276 23538 27328
rect 23566 27276 23572 27328
rect 23624 27316 23630 27328
rect 23753 27319 23811 27325
rect 23753 27316 23765 27319
rect 23624 27288 23765 27316
rect 23624 27276 23630 27288
rect 23753 27285 23765 27288
rect 23799 27285 23811 27319
rect 24136 27316 24164 27424
rect 24394 27384 24400 27396
rect 24355 27356 24400 27384
rect 24394 27344 24400 27356
rect 24452 27344 24458 27396
rect 24504 27384 24532 27424
rect 25777 27421 25789 27455
rect 25823 27421 25835 27455
rect 25777 27415 25835 27421
rect 25866 27412 25872 27464
rect 25924 27452 25930 27464
rect 26142 27452 26148 27464
rect 25924 27424 25969 27452
rect 26103 27424 26148 27452
rect 25924 27412 25930 27424
rect 26142 27412 26148 27424
rect 26200 27412 26206 27464
rect 26234 27412 26240 27464
rect 26292 27461 26298 27464
rect 26292 27452 26300 27461
rect 26292 27424 26337 27452
rect 26292 27415 26300 27424
rect 26292 27412 26298 27415
rect 26418 27412 26424 27464
rect 26476 27452 26482 27464
rect 27065 27455 27123 27461
rect 27065 27452 27077 27455
rect 26476 27424 27077 27452
rect 26476 27412 26482 27424
rect 27065 27421 27077 27424
rect 27111 27421 27123 27455
rect 27586 27452 27614 27492
rect 28184 27492 28540 27520
rect 27798 27452 27804 27464
rect 27586 27424 27804 27452
rect 27065 27415 27123 27421
rect 27798 27412 27804 27424
rect 27856 27412 27862 27464
rect 27949 27455 28007 27461
rect 27949 27421 27961 27455
rect 27995 27452 28007 27455
rect 28184 27452 28212 27492
rect 28534 27480 28540 27492
rect 28592 27480 28598 27532
rect 27995 27424 28212 27452
rect 27995 27421 28007 27424
rect 27949 27415 28007 27421
rect 28258 27412 28264 27464
rect 28316 27461 28322 27464
rect 28316 27452 28324 27461
rect 28316 27424 28361 27452
rect 28316 27415 28324 27424
rect 28316 27412 28322 27415
rect 26053 27387 26111 27393
rect 24504 27356 26004 27384
rect 24857 27319 24915 27325
rect 24857 27316 24869 27319
rect 24136 27288 24869 27316
rect 23753 27279 23811 27285
rect 24857 27285 24869 27288
rect 24903 27285 24915 27319
rect 25976 27316 26004 27356
rect 26053 27353 26065 27387
rect 26099 27384 26111 27387
rect 26510 27384 26516 27396
rect 26099 27356 26516 27384
rect 26099 27353 26111 27356
rect 26053 27347 26111 27353
rect 26510 27344 26516 27356
rect 26568 27344 26574 27396
rect 26881 27387 26939 27393
rect 26881 27353 26893 27387
rect 26927 27384 26939 27387
rect 27706 27384 27712 27396
rect 26927 27356 27712 27384
rect 26927 27353 26939 27356
rect 26881 27347 26939 27353
rect 26896 27316 26924 27347
rect 27706 27344 27712 27356
rect 27764 27344 27770 27396
rect 28074 27384 28080 27396
rect 28035 27356 28080 27384
rect 28074 27344 28080 27356
rect 28132 27344 28138 27396
rect 28169 27387 28227 27393
rect 28169 27353 28181 27387
rect 28215 27384 28227 27387
rect 28626 27384 28632 27396
rect 28215 27356 28632 27384
rect 28215 27353 28227 27356
rect 28169 27347 28227 27353
rect 28626 27344 28632 27356
rect 28684 27344 28690 27396
rect 29380 27384 29408 27560
rect 29914 27548 29920 27600
rect 29972 27548 29978 27600
rect 29730 27480 29736 27532
rect 29788 27520 29794 27532
rect 29932 27520 29960 27548
rect 29788 27492 29960 27520
rect 29788 27480 29794 27492
rect 29454 27412 29460 27464
rect 29512 27452 29518 27464
rect 29932 27461 29960 27492
rect 29825 27455 29883 27461
rect 29825 27452 29837 27455
rect 29512 27424 29837 27452
rect 29512 27412 29518 27424
rect 29825 27421 29837 27424
rect 29871 27421 29883 27455
rect 29825 27415 29883 27421
rect 29917 27455 29975 27461
rect 29917 27421 29929 27455
rect 29963 27421 29975 27455
rect 29917 27415 29975 27421
rect 30006 27412 30012 27464
rect 30064 27452 30070 27464
rect 30208 27461 30236 27616
rect 30193 27455 30251 27461
rect 30064 27424 30109 27452
rect 30064 27412 30070 27424
rect 30193 27421 30205 27455
rect 30239 27421 30251 27455
rect 30193 27415 30251 27421
rect 31386 27384 31392 27396
rect 29380 27356 31392 27384
rect 31386 27344 31392 27356
rect 31444 27344 31450 27396
rect 27246 27316 27252 27328
rect 25976 27288 26924 27316
rect 27207 27288 27252 27316
rect 24857 27279 24915 27285
rect 27246 27276 27252 27288
rect 27304 27276 27310 27328
rect 28445 27319 28503 27325
rect 28445 27285 28457 27319
rect 28491 27316 28503 27319
rect 28534 27316 28540 27328
rect 28491 27288 28540 27316
rect 28491 27285 28503 27288
rect 28445 27279 28503 27285
rect 28534 27276 28540 27288
rect 28592 27276 28598 27328
rect 29546 27316 29552 27328
rect 29507 27288 29552 27316
rect 29546 27276 29552 27288
rect 29604 27276 29610 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 6914 27112 6920 27124
rect 6380 27084 6920 27112
rect 5534 27044 5540 27056
rect 4448 27016 5540 27044
rect 4448 26985 4476 27016
rect 5534 27004 5540 27016
rect 5592 27004 5598 27056
rect 6380 27053 6408 27084
rect 6914 27072 6920 27084
rect 6972 27112 6978 27124
rect 7193 27115 7251 27121
rect 7193 27112 7205 27115
rect 6972 27084 7205 27112
rect 6972 27072 6978 27084
rect 7193 27081 7205 27084
rect 7239 27112 7251 27115
rect 7742 27112 7748 27124
rect 7239 27084 7748 27112
rect 7239 27081 7251 27084
rect 7193 27075 7251 27081
rect 7742 27072 7748 27084
rect 7800 27072 7806 27124
rect 7837 27115 7895 27121
rect 7837 27081 7849 27115
rect 7883 27112 7895 27115
rect 9214 27112 9220 27124
rect 7883 27084 9220 27112
rect 7883 27081 7895 27084
rect 7837 27075 7895 27081
rect 9214 27072 9220 27084
rect 9272 27072 9278 27124
rect 10410 27112 10416 27124
rect 10371 27084 10416 27112
rect 10410 27072 10416 27084
rect 10468 27072 10474 27124
rect 14274 27072 14280 27124
rect 14332 27112 14338 27124
rect 15286 27112 15292 27124
rect 14332 27084 15292 27112
rect 14332 27072 14338 27084
rect 15286 27072 15292 27084
rect 15344 27072 15350 27124
rect 15381 27115 15439 27121
rect 15381 27081 15393 27115
rect 15427 27112 15439 27115
rect 15470 27112 15476 27124
rect 15427 27084 15476 27112
rect 15427 27081 15439 27084
rect 15381 27075 15439 27081
rect 15470 27072 15476 27084
rect 15528 27072 15534 27124
rect 16758 27112 16764 27124
rect 15580 27084 16764 27112
rect 6365 27047 6423 27053
rect 6365 27013 6377 27047
rect 6411 27013 6423 27047
rect 6365 27007 6423 27013
rect 6454 27004 6460 27056
rect 6512 27044 6518 27056
rect 6565 27047 6623 27053
rect 6565 27044 6577 27047
rect 6512 27016 6577 27044
rect 6512 27004 6518 27016
rect 6565 27013 6577 27016
rect 6611 27013 6623 27047
rect 6565 27007 6623 27013
rect 4433 26979 4491 26985
rect 4433 26945 4445 26979
rect 4479 26945 4491 26979
rect 4433 26939 4491 26945
rect 4700 26979 4758 26985
rect 4700 26945 4712 26979
rect 4746 26976 4758 26979
rect 5442 26976 5448 26988
rect 4746 26948 5448 26976
rect 4746 26945 4758 26948
rect 4700 26939 4758 26945
rect 5442 26936 5448 26948
rect 5500 26936 5506 26988
rect 7190 26936 7196 26988
rect 7248 26976 7254 26988
rect 7377 26979 7435 26985
rect 7377 26976 7389 26979
rect 7248 26948 7389 26976
rect 7248 26936 7254 26948
rect 7377 26945 7389 26948
rect 7423 26945 7435 26979
rect 7377 26939 7435 26945
rect 8021 26979 8079 26985
rect 8021 26945 8033 26979
rect 8067 26976 8079 26979
rect 8110 26976 8116 26988
rect 8067 26948 8116 26976
rect 8067 26945 8079 26948
rect 8021 26939 8079 26945
rect 8110 26936 8116 26948
rect 8168 26936 8174 26988
rect 8662 26976 8668 26988
rect 8623 26948 8668 26976
rect 8662 26936 8668 26948
rect 8720 26936 8726 26988
rect 9950 26976 9956 26988
rect 9911 26948 9956 26976
rect 9950 26936 9956 26948
rect 10008 26936 10014 26988
rect 10594 26976 10600 26988
rect 10555 26948 10600 26976
rect 10594 26936 10600 26948
rect 10652 26936 10658 26988
rect 13909 26979 13967 26985
rect 13909 26945 13921 26979
rect 13955 26976 13967 26979
rect 14366 26976 14372 26988
rect 13955 26948 14372 26976
rect 13955 26945 13967 26948
rect 13909 26939 13967 26945
rect 14366 26936 14372 26948
rect 14424 26976 14430 26988
rect 14734 26976 14740 26988
rect 14424 26948 14740 26976
rect 14424 26936 14430 26948
rect 14734 26936 14740 26948
rect 14792 26936 14798 26988
rect 15580 26976 15608 27084
rect 16758 27072 16764 27084
rect 16816 27072 16822 27124
rect 17218 27112 17224 27124
rect 17179 27084 17224 27112
rect 17218 27072 17224 27084
rect 17276 27112 17282 27124
rect 17276 27084 23152 27112
rect 17276 27072 17282 27084
rect 19426 27044 19432 27056
rect 18616 27016 19432 27044
rect 15657 26979 15715 26985
rect 15657 26976 15669 26979
rect 15580 26948 15669 26976
rect 15657 26945 15669 26948
rect 15703 26945 15715 26979
rect 15657 26939 15715 26945
rect 15749 26979 15807 26985
rect 15749 26945 15761 26979
rect 15795 26945 15807 26979
rect 15749 26939 15807 26945
rect 13170 26868 13176 26920
rect 13228 26908 13234 26920
rect 13541 26911 13599 26917
rect 13541 26908 13553 26911
rect 13228 26880 13553 26908
rect 13228 26868 13234 26880
rect 13541 26877 13553 26880
rect 13587 26877 13599 26911
rect 13541 26871 13599 26877
rect 13814 26868 13820 26920
rect 13872 26908 13878 26920
rect 14001 26911 14059 26917
rect 14001 26908 14013 26911
rect 13872 26880 14013 26908
rect 13872 26868 13878 26880
rect 14001 26877 14013 26880
rect 14047 26908 14059 26911
rect 15102 26908 15108 26920
rect 14047 26880 15108 26908
rect 14047 26877 14059 26880
rect 14001 26871 14059 26877
rect 15102 26868 15108 26880
rect 15160 26868 15166 26920
rect 5813 26775 5871 26781
rect 5813 26741 5825 26775
rect 5859 26772 5871 26775
rect 6549 26775 6607 26781
rect 6549 26772 6561 26775
rect 5859 26744 6561 26772
rect 5859 26741 5871 26744
rect 5813 26735 5871 26741
rect 6549 26741 6561 26744
rect 6595 26741 6607 26775
rect 6730 26772 6736 26784
rect 6691 26744 6736 26772
rect 6549 26735 6607 26741
rect 6730 26732 6736 26744
rect 6788 26732 6794 26784
rect 8478 26772 8484 26784
rect 8439 26744 8484 26772
rect 8478 26732 8484 26744
rect 8536 26732 8542 26784
rect 9766 26772 9772 26784
rect 9727 26744 9772 26772
rect 9766 26732 9772 26744
rect 9824 26732 9830 26784
rect 14185 26775 14243 26781
rect 14185 26741 14197 26775
rect 14231 26772 14243 26775
rect 14274 26772 14280 26784
rect 14231 26744 14280 26772
rect 14231 26741 14243 26744
rect 14185 26735 14243 26741
rect 14274 26732 14280 26744
rect 14332 26732 14338 26784
rect 15764 26772 15792 26939
rect 15838 26936 15844 26988
rect 15896 26976 15902 26988
rect 16025 26979 16083 26985
rect 15896 26948 15941 26976
rect 15896 26936 15902 26948
rect 16025 26945 16037 26979
rect 16071 26945 16083 26979
rect 16025 26939 16083 26945
rect 17129 26979 17187 26985
rect 17129 26945 17141 26979
rect 17175 26945 17187 26979
rect 17954 26976 17960 26988
rect 17915 26948 17960 26976
rect 17129 26939 17187 26945
rect 16040 26840 16068 26939
rect 17144 26908 17172 26939
rect 17954 26936 17960 26948
rect 18012 26936 18018 26988
rect 18616 26985 18644 27016
rect 19426 27004 19432 27016
rect 19484 27044 19490 27056
rect 20622 27044 20628 27056
rect 19484 27016 20628 27044
rect 19484 27004 19490 27016
rect 20622 27004 20628 27016
rect 20680 27004 20686 27056
rect 22465 27047 22523 27053
rect 22465 27044 22477 27047
rect 21008 27016 22477 27044
rect 18601 26979 18659 26985
rect 18601 26945 18613 26979
rect 18647 26945 18659 26979
rect 18601 26939 18659 26945
rect 18690 26936 18696 26988
rect 18748 26936 18754 26988
rect 18868 26979 18926 26985
rect 18868 26945 18880 26979
rect 18914 26976 18926 26979
rect 19242 26976 19248 26988
rect 18914 26948 19248 26976
rect 18914 26945 18926 26948
rect 18868 26939 18926 26945
rect 19242 26936 19248 26948
rect 19300 26936 19306 26988
rect 19978 26936 19984 26988
rect 20036 26976 20042 26988
rect 21008 26985 21036 27016
rect 22465 27013 22477 27016
rect 22511 27013 22523 27047
rect 23124 27044 23152 27084
rect 23842 27072 23848 27124
rect 23900 27112 23906 27124
rect 24121 27115 24179 27121
rect 24121 27112 24133 27115
rect 23900 27084 24133 27112
rect 23900 27072 23906 27084
rect 24121 27081 24133 27084
rect 24167 27081 24179 27115
rect 24121 27075 24179 27081
rect 24210 27072 24216 27124
rect 24268 27112 24274 27124
rect 24765 27115 24823 27121
rect 24765 27112 24777 27115
rect 24268 27084 24777 27112
rect 24268 27072 24274 27084
rect 24765 27081 24777 27084
rect 24811 27081 24823 27115
rect 24765 27075 24823 27081
rect 25314 27072 25320 27124
rect 25372 27112 25378 27124
rect 25409 27115 25467 27121
rect 25409 27112 25421 27115
rect 25372 27084 25421 27112
rect 25372 27072 25378 27084
rect 25409 27081 25421 27084
rect 25455 27081 25467 27115
rect 25866 27112 25872 27124
rect 25409 27075 25467 27081
rect 25792 27084 25872 27112
rect 23198 27044 23204 27056
rect 23111 27016 23204 27044
rect 22465 27007 22523 27013
rect 23198 27004 23204 27016
rect 23256 27004 23262 27056
rect 25792 27044 25820 27084
rect 25866 27072 25872 27084
rect 25924 27072 25930 27124
rect 28077 27115 28135 27121
rect 28077 27081 28089 27115
rect 28123 27112 28135 27115
rect 28994 27112 29000 27124
rect 28123 27084 29000 27112
rect 28123 27081 28135 27084
rect 28077 27075 28135 27081
rect 28994 27072 29000 27084
rect 29052 27072 29058 27124
rect 29086 27072 29092 27124
rect 29144 27112 29150 27124
rect 31205 27115 31263 27121
rect 31205 27112 31217 27115
rect 29144 27084 31217 27112
rect 29144 27072 29150 27084
rect 31205 27081 31217 27084
rect 31251 27081 31263 27115
rect 31205 27075 31263 27081
rect 27246 27044 27252 27056
rect 24044 27016 25820 27044
rect 25884 27016 27252 27044
rect 24044 26988 24072 27016
rect 20993 26979 21051 26985
rect 20036 26948 20944 26976
rect 20036 26936 20042 26948
rect 18141 26911 18199 26917
rect 18141 26908 18153 26911
rect 17144 26880 18153 26908
rect 18141 26877 18153 26880
rect 18187 26908 18199 26911
rect 18708 26908 18736 26936
rect 20806 26908 20812 26920
rect 18187 26880 18736 26908
rect 19996 26880 20812 26908
rect 18187 26877 18199 26880
rect 18141 26871 18199 26877
rect 19996 26852 20024 26880
rect 20806 26868 20812 26880
rect 20864 26868 20870 26920
rect 19978 26840 19984 26852
rect 16040 26812 17816 26840
rect 19891 26812 19984 26840
rect 17788 26784 17816 26812
rect 19978 26800 19984 26812
rect 20036 26800 20042 26852
rect 20916 26840 20944 26948
rect 20993 26945 21005 26979
rect 21039 26945 21051 26979
rect 20993 26939 21051 26945
rect 21177 26979 21235 26985
rect 21177 26945 21189 26979
rect 21223 26945 21235 26979
rect 21177 26939 21235 26945
rect 21192 26908 21220 26939
rect 21266 26936 21272 26988
rect 21324 26976 21330 26988
rect 22278 26976 22284 26988
rect 21324 26948 21369 26976
rect 22239 26948 22284 26976
rect 21324 26936 21330 26948
rect 22278 26936 22284 26948
rect 22336 26936 22342 26988
rect 22830 26936 22836 26988
rect 22888 26936 22894 26988
rect 23385 26979 23443 26985
rect 23385 26945 23397 26979
rect 23431 26945 23443 26979
rect 24026 26976 24032 26988
rect 23987 26948 24032 26976
rect 23385 26939 23443 26945
rect 21726 26908 21732 26920
rect 21192 26880 21732 26908
rect 21726 26868 21732 26880
rect 21784 26868 21790 26920
rect 21821 26911 21879 26917
rect 21821 26877 21833 26911
rect 21867 26877 21879 26911
rect 21821 26871 21879 26877
rect 22189 26911 22247 26917
rect 22189 26877 22201 26911
rect 22235 26908 22247 26911
rect 22848 26908 22876 26936
rect 22235 26880 22876 26908
rect 23400 26908 23428 26939
rect 24026 26936 24032 26948
rect 24084 26936 24090 26988
rect 24210 26976 24216 26988
rect 24171 26948 24216 26976
rect 24210 26936 24216 26948
rect 24268 26936 24274 26988
rect 24688 26985 24716 27016
rect 24673 26979 24731 26985
rect 24673 26945 24685 26979
rect 24719 26945 24731 26979
rect 24673 26939 24731 26945
rect 24857 26979 24915 26985
rect 24857 26945 24869 26979
rect 24903 26945 24915 26979
rect 24857 26939 24915 26945
rect 24228 26908 24256 26936
rect 24872 26908 24900 26939
rect 25590 26936 25596 26988
rect 25648 26976 25654 26988
rect 25884 26985 25912 27016
rect 27246 27004 27252 27016
rect 27304 27004 27310 27056
rect 27706 27044 27712 27056
rect 27667 27016 27712 27044
rect 27706 27004 27712 27016
rect 27764 27004 27770 27056
rect 27816 27016 28120 27044
rect 25685 26979 25743 26985
rect 25685 26976 25697 26979
rect 25648 26948 25697 26976
rect 25648 26936 25654 26948
rect 25685 26945 25697 26948
rect 25731 26945 25743 26979
rect 25685 26939 25743 26945
rect 25777 26979 25835 26985
rect 25777 26945 25789 26979
rect 25823 26945 25835 26979
rect 25777 26939 25835 26945
rect 25869 26979 25927 26985
rect 25869 26945 25881 26979
rect 25915 26945 25927 26979
rect 26053 26979 26111 26985
rect 26053 26976 26065 26979
rect 25869 26939 25927 26945
rect 25976 26948 26065 26976
rect 23400 26880 24900 26908
rect 22235 26877 22247 26880
rect 22189 26871 22247 26877
rect 21836 26840 21864 26871
rect 22296 26852 22324 26880
rect 25498 26868 25504 26920
rect 25556 26908 25562 26920
rect 25792 26908 25820 26939
rect 25556 26880 25820 26908
rect 25556 26868 25562 26880
rect 20916 26812 21864 26840
rect 22278 26800 22284 26852
rect 22336 26800 22342 26852
rect 23290 26800 23296 26852
rect 23348 26840 23354 26852
rect 25976 26840 26004 26948
rect 26053 26945 26065 26948
rect 26099 26976 26111 26979
rect 26786 26976 26792 26988
rect 26099 26948 26792 26976
rect 26099 26945 26111 26948
rect 26053 26939 26111 26945
rect 26786 26936 26792 26948
rect 26844 26936 26850 26988
rect 26970 26936 26976 26988
rect 27028 26976 27034 26988
rect 27065 26979 27123 26985
rect 27065 26976 27077 26979
rect 27028 26948 27077 26976
rect 27028 26936 27034 26948
rect 27065 26945 27077 26948
rect 27111 26976 27123 26979
rect 27816 26976 27844 27016
rect 27111 26948 27844 26976
rect 27111 26945 27123 26948
rect 27065 26939 27123 26945
rect 27890 26936 27896 26988
rect 27948 26976 27954 26988
rect 28092 26976 28120 27016
rect 28350 27004 28356 27056
rect 28408 27044 28414 27056
rect 28902 27044 28908 27056
rect 28408 27016 28580 27044
rect 28863 27016 28908 27044
rect 28408 27004 28414 27016
rect 28552 26985 28580 27016
rect 28902 27004 28908 27016
rect 28960 27004 28966 27056
rect 29546 27004 29552 27056
rect 29604 27044 29610 27056
rect 30070 27047 30128 27053
rect 30070 27044 30082 27047
rect 29604 27016 30082 27044
rect 29604 27004 29610 27016
rect 30070 27013 30082 27016
rect 30116 27013 30128 27047
rect 30070 27007 30128 27013
rect 28718 26985 28724 26988
rect 28537 26979 28595 26985
rect 27948 26948 27993 26976
rect 28092 26948 28488 26976
rect 27948 26936 27954 26948
rect 26510 26868 26516 26920
rect 26568 26908 26574 26920
rect 26988 26908 27016 26936
rect 26568 26880 27016 26908
rect 26568 26868 26574 26880
rect 27798 26868 27804 26920
rect 27856 26908 27862 26920
rect 28166 26908 28172 26920
rect 27856 26880 28172 26908
rect 27856 26868 27862 26880
rect 28166 26868 28172 26880
rect 28224 26868 28230 26920
rect 28460 26908 28488 26948
rect 28537 26945 28549 26979
rect 28583 26945 28595 26979
rect 28537 26939 28595 26945
rect 28685 26979 28724 26985
rect 28685 26945 28697 26979
rect 28685 26939 28724 26945
rect 28718 26936 28724 26939
rect 28776 26936 28782 26988
rect 28813 26979 28871 26985
rect 28813 26945 28825 26979
rect 28859 26945 28871 26979
rect 29002 26979 29060 26985
rect 29002 26976 29014 26979
rect 28813 26939 28871 26945
rect 28920 26948 29014 26976
rect 28828 26908 28856 26939
rect 28460 26880 28856 26908
rect 23348 26812 26004 26840
rect 27249 26843 27307 26849
rect 23348 26800 23354 26812
rect 27249 26809 27261 26843
rect 27295 26840 27307 26843
rect 28074 26840 28080 26852
rect 27295 26812 28080 26840
rect 27295 26809 27307 26812
rect 27249 26803 27307 26809
rect 28074 26800 28080 26812
rect 28132 26800 28138 26852
rect 16758 26772 16764 26784
rect 15764 26744 16764 26772
rect 16758 26732 16764 26744
rect 16816 26732 16822 26784
rect 17770 26732 17776 26784
rect 17828 26772 17834 26784
rect 20254 26772 20260 26784
rect 17828 26744 20260 26772
rect 17828 26732 17834 26744
rect 20254 26732 20260 26744
rect 20312 26732 20318 26784
rect 20809 26775 20867 26781
rect 20809 26741 20821 26775
rect 20855 26772 20867 26775
rect 20898 26772 20904 26784
rect 20855 26744 20904 26772
rect 20855 26741 20867 26744
rect 20809 26735 20867 26741
rect 20898 26732 20904 26744
rect 20956 26732 20962 26784
rect 23106 26732 23112 26784
rect 23164 26772 23170 26784
rect 23569 26775 23627 26781
rect 23569 26772 23581 26775
rect 23164 26744 23581 26772
rect 23164 26732 23170 26744
rect 23569 26741 23581 26744
rect 23615 26741 23627 26775
rect 23569 26735 23627 26741
rect 26234 26732 26240 26784
rect 26292 26772 26298 26784
rect 28920 26772 28948 26948
rect 29002 26945 29014 26948
rect 29048 26976 29060 26979
rect 29178 26976 29184 26988
rect 29048 26948 29184 26976
rect 29048 26945 29060 26948
rect 29002 26939 29060 26945
rect 29178 26936 29184 26948
rect 29236 26936 29242 26988
rect 29825 26911 29883 26917
rect 29825 26877 29837 26911
rect 29871 26877 29883 26911
rect 29825 26871 29883 26877
rect 26292 26744 28948 26772
rect 26292 26732 26298 26744
rect 29086 26732 29092 26784
rect 29144 26772 29150 26784
rect 29181 26775 29239 26781
rect 29181 26772 29193 26775
rect 29144 26744 29193 26772
rect 29144 26732 29150 26744
rect 29181 26741 29193 26744
rect 29227 26741 29239 26775
rect 29840 26772 29868 26871
rect 30098 26772 30104 26784
rect 29840 26744 30104 26772
rect 29181 26735 29239 26741
rect 30098 26732 30104 26744
rect 30156 26732 30162 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 11514 26568 11520 26580
rect 11256 26540 11520 26568
rect 11256 26441 11284 26540
rect 11514 26528 11520 26540
rect 11572 26528 11578 26580
rect 12621 26571 12679 26577
rect 12621 26537 12633 26571
rect 12667 26568 12679 26571
rect 12894 26568 12900 26580
rect 12667 26540 12900 26568
rect 12667 26537 12679 26540
rect 12621 26531 12679 26537
rect 12894 26528 12900 26540
rect 12952 26528 12958 26580
rect 14458 26528 14464 26580
rect 14516 26568 14522 26580
rect 15473 26571 15531 26577
rect 15473 26568 15485 26571
rect 14516 26540 15485 26568
rect 14516 26528 14522 26540
rect 15473 26537 15485 26540
rect 15519 26537 15531 26571
rect 26234 26568 26240 26580
rect 15473 26531 15531 26537
rect 15580 26540 26240 26568
rect 11241 26435 11299 26441
rect 11241 26401 11253 26435
rect 11287 26401 11299 26435
rect 12912 26432 12940 26528
rect 13262 26460 13268 26512
rect 13320 26500 13326 26512
rect 15580 26500 15608 26540
rect 26234 26528 26240 26540
rect 26292 26528 26298 26580
rect 28813 26571 28871 26577
rect 28813 26537 28825 26571
rect 28859 26568 28871 26571
rect 30006 26568 30012 26580
rect 28859 26540 30012 26568
rect 28859 26537 28871 26540
rect 28813 26531 28871 26537
rect 30006 26528 30012 26540
rect 30064 26528 30070 26580
rect 31386 26568 31392 26580
rect 31347 26540 31392 26568
rect 31386 26528 31392 26540
rect 31444 26528 31450 26580
rect 13320 26472 13584 26500
rect 13320 26460 13326 26472
rect 13556 26432 13584 26472
rect 15120 26472 15608 26500
rect 12912 26404 13492 26432
rect 13556 26404 14228 26432
rect 11241 26395 11299 26401
rect 4893 26367 4951 26373
rect 4893 26333 4905 26367
rect 4939 26364 4951 26367
rect 5534 26364 5540 26376
rect 4939 26336 5540 26364
rect 4939 26333 4951 26336
rect 4893 26327 4951 26333
rect 5534 26324 5540 26336
rect 5592 26324 5598 26376
rect 7009 26367 7067 26373
rect 7009 26333 7021 26367
rect 7055 26364 7067 26367
rect 8941 26367 8999 26373
rect 8941 26364 8953 26367
rect 7055 26336 8953 26364
rect 7055 26333 7067 26336
rect 7009 26327 7067 26333
rect 8941 26333 8953 26336
rect 8987 26364 8999 26367
rect 9030 26364 9036 26376
rect 8987 26336 9036 26364
rect 8987 26333 8999 26336
rect 8941 26327 8999 26333
rect 9030 26324 9036 26336
rect 9088 26324 9094 26376
rect 13262 26364 13268 26376
rect 13223 26336 13268 26364
rect 13262 26324 13268 26336
rect 13320 26324 13326 26376
rect 13464 26373 13492 26404
rect 13449 26367 13507 26373
rect 13449 26333 13461 26367
rect 13495 26333 13507 26367
rect 13449 26327 13507 26333
rect 13541 26367 13599 26373
rect 13541 26333 13553 26367
rect 13587 26333 13599 26367
rect 14090 26364 14096 26376
rect 14051 26336 14096 26364
rect 13541 26327 13599 26333
rect 5160 26299 5218 26305
rect 5160 26265 5172 26299
rect 5206 26296 5218 26299
rect 5626 26296 5632 26308
rect 5206 26268 5632 26296
rect 5206 26265 5218 26268
rect 5160 26259 5218 26265
rect 5626 26256 5632 26268
rect 5684 26256 5690 26308
rect 7276 26299 7334 26305
rect 7276 26265 7288 26299
rect 7322 26296 7334 26299
rect 8478 26296 8484 26308
rect 7322 26268 8484 26296
rect 7322 26265 7334 26268
rect 7276 26259 7334 26265
rect 8478 26256 8484 26268
rect 8536 26256 8542 26308
rect 9208 26299 9266 26305
rect 9208 26265 9220 26299
rect 9254 26296 9266 26299
rect 10778 26296 10784 26308
rect 9254 26268 10784 26296
rect 9254 26265 9266 26268
rect 9208 26259 9266 26265
rect 10778 26256 10784 26268
rect 10836 26256 10842 26308
rect 11508 26299 11566 26305
rect 11508 26265 11520 26299
rect 11554 26296 11566 26299
rect 13081 26299 13139 26305
rect 13081 26296 13093 26299
rect 11554 26268 13093 26296
rect 11554 26265 11566 26268
rect 11508 26259 11566 26265
rect 13081 26265 13093 26268
rect 13127 26265 13139 26299
rect 13556 26296 13584 26327
rect 14090 26324 14096 26336
rect 14148 26324 14154 26376
rect 14200 26364 14228 26404
rect 15120 26364 15148 26472
rect 21726 26460 21732 26512
rect 21784 26500 21790 26512
rect 22005 26503 22063 26509
rect 22005 26500 22017 26503
rect 21784 26472 22017 26500
rect 21784 26460 21790 26472
rect 22005 26469 22017 26472
rect 22051 26500 22063 26503
rect 24026 26500 24032 26512
rect 22051 26472 24032 26500
rect 22051 26469 22063 26472
rect 22005 26463 22063 26469
rect 24026 26460 24032 26472
rect 24084 26460 24090 26512
rect 15194 26392 15200 26444
rect 15252 26432 15258 26444
rect 18966 26432 18972 26444
rect 15252 26404 18972 26432
rect 15252 26392 15258 26404
rect 18966 26392 18972 26404
rect 19024 26432 19030 26444
rect 19521 26435 19579 26441
rect 19521 26432 19533 26435
rect 19024 26404 19533 26432
rect 19024 26392 19030 26404
rect 19521 26401 19533 26404
rect 19567 26401 19579 26435
rect 20622 26432 20628 26444
rect 20583 26404 20628 26432
rect 19521 26395 19579 26401
rect 20622 26392 20628 26404
rect 20680 26392 20686 26444
rect 23750 26432 23756 26444
rect 22940 26404 23756 26432
rect 22940 26376 22968 26404
rect 23750 26392 23756 26404
rect 23808 26392 23814 26444
rect 14200 26336 15148 26364
rect 17954 26324 17960 26376
rect 18012 26364 18018 26376
rect 18690 26364 18696 26376
rect 18012 26336 18696 26364
rect 18012 26324 18018 26336
rect 18690 26324 18696 26336
rect 18748 26364 18754 26376
rect 20898 26373 20904 26376
rect 19245 26367 19303 26373
rect 19245 26364 19257 26367
rect 18748 26336 19257 26364
rect 18748 26324 18754 26336
rect 19245 26333 19257 26336
rect 19291 26333 19303 26367
rect 20892 26364 20904 26373
rect 20859 26336 20904 26364
rect 19245 26327 19303 26333
rect 20892 26327 20904 26336
rect 20898 26324 20904 26327
rect 20956 26324 20962 26376
rect 22922 26364 22928 26376
rect 22883 26336 22928 26364
rect 22922 26324 22928 26336
rect 22980 26324 22986 26376
rect 23017 26367 23075 26373
rect 23017 26333 23029 26367
rect 23063 26333 23075 26367
rect 23017 26327 23075 26333
rect 13556 26268 14136 26296
rect 13081 26259 13139 26265
rect 6273 26231 6331 26237
rect 6273 26197 6285 26231
rect 6319 26228 6331 26231
rect 6546 26228 6552 26240
rect 6319 26200 6552 26228
rect 6319 26197 6331 26200
rect 6273 26191 6331 26197
rect 6546 26188 6552 26200
rect 6604 26188 6610 26240
rect 8386 26228 8392 26240
rect 8347 26200 8392 26228
rect 8386 26188 8392 26200
rect 8444 26188 8450 26240
rect 10042 26188 10048 26240
rect 10100 26228 10106 26240
rect 10321 26231 10379 26237
rect 10321 26228 10333 26231
rect 10100 26200 10333 26228
rect 10100 26188 10106 26200
rect 10321 26197 10333 26200
rect 10367 26197 10379 26231
rect 14108 26228 14136 26268
rect 14182 26256 14188 26308
rect 14240 26296 14246 26308
rect 14338 26299 14396 26305
rect 14338 26296 14350 26299
rect 14240 26268 14350 26296
rect 14240 26256 14246 26268
rect 14338 26265 14350 26268
rect 14384 26265 14396 26299
rect 14338 26259 14396 26265
rect 15286 26256 15292 26308
rect 15344 26296 15350 26308
rect 23032 26296 23060 26327
rect 23106 26324 23112 26376
rect 23164 26364 23170 26376
rect 23164 26336 23209 26364
rect 23164 26324 23170 26336
rect 23290 26324 23296 26376
rect 23348 26364 23354 26376
rect 23348 26336 23393 26364
rect 23348 26324 23354 26336
rect 27706 26324 27712 26376
rect 27764 26364 27770 26376
rect 28445 26367 28503 26373
rect 28445 26364 28457 26367
rect 27764 26336 28457 26364
rect 27764 26324 27770 26336
rect 28445 26333 28457 26336
rect 28491 26333 28503 26367
rect 28445 26327 28503 26333
rect 28629 26367 28687 26373
rect 28629 26333 28641 26367
rect 28675 26364 28687 26367
rect 28994 26364 29000 26376
rect 28675 26336 29000 26364
rect 28675 26333 28687 26336
rect 28629 26327 28687 26333
rect 28994 26324 29000 26336
rect 29052 26324 29058 26376
rect 30009 26367 30067 26373
rect 30009 26333 30021 26367
rect 30055 26364 30067 26367
rect 30098 26364 30104 26376
rect 30055 26336 30104 26364
rect 30055 26333 30067 26336
rect 30009 26327 30067 26333
rect 30098 26324 30104 26336
rect 30156 26324 30162 26376
rect 30282 26373 30288 26376
rect 30276 26364 30288 26373
rect 30243 26336 30288 26364
rect 30276 26327 30288 26336
rect 30282 26324 30288 26327
rect 30340 26324 30346 26376
rect 25498 26296 25504 26308
rect 15344 26268 25504 26296
rect 15344 26256 15350 26268
rect 25498 26256 25504 26268
rect 25556 26296 25562 26308
rect 29730 26296 29736 26308
rect 25556 26268 29736 26296
rect 25556 26256 25562 26268
rect 29730 26256 29736 26268
rect 29788 26256 29794 26308
rect 14642 26228 14648 26240
rect 14108 26200 14648 26228
rect 10321 26191 10379 26197
rect 14642 26188 14648 26200
rect 14700 26188 14706 26240
rect 22649 26231 22707 26237
rect 22649 26197 22661 26231
rect 22695 26228 22707 26231
rect 22738 26228 22744 26240
rect 22695 26200 22744 26228
rect 22695 26197 22707 26200
rect 22649 26191 22707 26197
rect 22738 26188 22744 26200
rect 22796 26188 22802 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 5537 26027 5595 26033
rect 5537 25993 5549 26027
rect 5583 26024 5595 26027
rect 5626 26024 5632 26036
rect 5583 25996 5632 26024
rect 5583 25993 5595 25996
rect 5537 25987 5595 25993
rect 5626 25984 5632 25996
rect 5684 25984 5690 26036
rect 6914 26024 6920 26036
rect 6380 25996 6920 26024
rect 6380 25965 6408 25996
rect 6914 25984 6920 25996
rect 6972 26024 6978 26036
rect 8113 26027 8171 26033
rect 6972 25996 7788 26024
rect 6972 25984 6978 25996
rect 6365 25959 6423 25965
rect 6365 25925 6377 25959
rect 6411 25925 6423 25959
rect 6365 25919 6423 25925
rect 6454 25916 6460 25968
rect 6512 25956 6518 25968
rect 7760 25965 7788 25996
rect 8113 25993 8125 26027
rect 8159 26024 8171 26027
rect 8662 26024 8668 26036
rect 8159 25996 8668 26024
rect 8159 25993 8171 25996
rect 8113 25987 8171 25993
rect 8662 25984 8668 25996
rect 8720 25984 8726 26036
rect 10778 26024 10784 26036
rect 10739 25996 10784 26024
rect 10778 25984 10784 25996
rect 10836 25984 10842 26036
rect 13262 25984 13268 26036
rect 13320 26024 13326 26036
rect 13633 26027 13691 26033
rect 13633 26024 13645 26027
rect 13320 25996 13645 26024
rect 13320 25984 13326 25996
rect 13633 25993 13645 25996
rect 13679 25993 13691 26027
rect 13633 25987 13691 25993
rect 14093 26027 14151 26033
rect 14093 25993 14105 26027
rect 14139 26024 14151 26027
rect 14182 26024 14188 26036
rect 14139 25996 14188 26024
rect 14139 25993 14151 25996
rect 14093 25987 14151 25993
rect 14182 25984 14188 25996
rect 14240 25984 14246 26036
rect 14458 26024 14464 26036
rect 14419 25996 14464 26024
rect 14458 25984 14464 25996
rect 14516 25984 14522 26036
rect 15933 26027 15991 26033
rect 15933 25993 15945 26027
rect 15979 26024 15991 26027
rect 16298 26024 16304 26036
rect 15979 25996 16304 26024
rect 15979 25993 15991 25996
rect 15933 25987 15991 25993
rect 16298 25984 16304 25996
rect 16356 25984 16362 26036
rect 16942 26024 16948 26036
rect 16776 25996 16948 26024
rect 6565 25959 6623 25965
rect 6565 25956 6577 25959
rect 6512 25928 6577 25956
rect 6512 25916 6518 25928
rect 6565 25925 6577 25928
rect 6611 25956 6623 25959
rect 7745 25959 7803 25965
rect 6611 25928 7696 25956
rect 6611 25925 6623 25928
rect 6565 25919 6623 25925
rect 5721 25891 5779 25897
rect 5721 25857 5733 25891
rect 5767 25888 5779 25891
rect 7668 25888 7696 25928
rect 7745 25925 7757 25959
rect 7791 25925 7803 25959
rect 7945 25959 8003 25965
rect 7945 25956 7957 25959
rect 7745 25919 7803 25925
rect 7944 25925 7957 25956
rect 7991 25956 8003 25959
rect 9766 25956 9772 25968
rect 7991 25928 9772 25956
rect 7991 25925 8003 25928
rect 7944 25919 8003 25925
rect 7944 25888 7972 25919
rect 9766 25916 9772 25928
rect 9824 25916 9830 25968
rect 15565 25959 15623 25965
rect 15565 25925 15577 25959
rect 15611 25956 15623 25959
rect 16666 25956 16672 25968
rect 15611 25928 16672 25956
rect 15611 25925 15623 25928
rect 15565 25919 15623 25925
rect 16666 25916 16672 25928
rect 16724 25916 16730 25968
rect 5767 25860 6776 25888
rect 7668 25860 7972 25888
rect 8941 25891 8999 25897
rect 5767 25857 5779 25860
rect 5721 25851 5779 25857
rect 6748 25761 6776 25860
rect 8941 25857 8953 25891
rect 8987 25888 8999 25891
rect 9030 25888 9036 25900
rect 8987 25860 9036 25888
rect 8987 25857 8999 25860
rect 8941 25851 8999 25857
rect 9030 25848 9036 25860
rect 9088 25848 9094 25900
rect 9208 25891 9266 25897
rect 9208 25857 9220 25891
rect 9254 25888 9266 25891
rect 9582 25888 9588 25900
rect 9254 25860 9588 25888
rect 9254 25857 9266 25860
rect 9208 25851 9266 25857
rect 9582 25848 9588 25860
rect 9640 25848 9646 25900
rect 10226 25848 10232 25900
rect 10284 25888 10290 25900
rect 10965 25891 11023 25897
rect 10965 25888 10977 25891
rect 10284 25860 10977 25888
rect 10284 25848 10290 25860
rect 10965 25857 10977 25860
rect 11011 25857 11023 25891
rect 10965 25851 11023 25857
rect 13449 25891 13507 25897
rect 13449 25857 13461 25891
rect 13495 25888 13507 25891
rect 13814 25888 13820 25900
rect 13495 25860 13820 25888
rect 13495 25857 13507 25860
rect 13449 25851 13507 25857
rect 13814 25848 13820 25860
rect 13872 25848 13878 25900
rect 14274 25888 14280 25900
rect 14235 25860 14280 25888
rect 14274 25848 14280 25860
rect 14332 25848 14338 25900
rect 14553 25891 14611 25897
rect 14553 25857 14565 25891
rect 14599 25888 14611 25891
rect 14642 25888 14648 25900
rect 14599 25860 14648 25888
rect 14599 25857 14611 25860
rect 14553 25851 14611 25857
rect 14642 25848 14648 25860
rect 14700 25848 14706 25900
rect 15286 25848 15292 25900
rect 15344 25888 15350 25900
rect 15749 25891 15807 25897
rect 15749 25888 15761 25891
rect 15344 25860 15761 25888
rect 15344 25848 15350 25860
rect 15749 25857 15761 25860
rect 15795 25888 15807 25891
rect 16776 25888 16804 25996
rect 16942 25984 16948 25996
rect 17000 25984 17006 26036
rect 18233 26027 18291 26033
rect 18233 25993 18245 26027
rect 18279 26024 18291 26027
rect 18414 26024 18420 26036
rect 18279 25996 18420 26024
rect 18279 25993 18291 25996
rect 18233 25987 18291 25993
rect 18414 25984 18420 25996
rect 18472 25984 18478 26036
rect 19334 26024 19340 26036
rect 19295 25996 19340 26024
rect 19334 25984 19340 25996
rect 19392 25984 19398 26036
rect 21085 26027 21143 26033
rect 21085 25993 21097 26027
rect 21131 26024 21143 26027
rect 21266 26024 21272 26036
rect 21131 25996 21272 26024
rect 21131 25993 21143 25996
rect 21085 25987 21143 25993
rect 21266 25984 21272 25996
rect 21324 25984 21330 26036
rect 24854 25984 24860 26036
rect 24912 26024 24918 26036
rect 25225 26027 25283 26033
rect 25225 26024 25237 26027
rect 24912 25996 25237 26024
rect 24912 25984 24918 25996
rect 25225 25993 25237 25996
rect 25271 25993 25283 26027
rect 26234 26024 26240 26036
rect 25225 25987 25283 25993
rect 25792 25996 26240 26024
rect 17310 25956 17316 25968
rect 16868 25928 17316 25956
rect 16868 25897 16896 25928
rect 17310 25916 17316 25928
rect 17368 25916 17374 25968
rect 18966 25956 18972 25968
rect 18927 25928 18972 25956
rect 18966 25916 18972 25928
rect 19024 25916 19030 25968
rect 19153 25959 19211 25965
rect 19153 25925 19165 25959
rect 19199 25956 19211 25959
rect 19978 25956 19984 25968
rect 19199 25928 19984 25956
rect 19199 25925 19211 25928
rect 19153 25919 19211 25925
rect 19978 25916 19984 25928
rect 20036 25916 20042 25968
rect 20257 25959 20315 25965
rect 20257 25925 20269 25959
rect 20303 25956 20315 25959
rect 20303 25928 21588 25956
rect 20303 25925 20315 25928
rect 20257 25919 20315 25925
rect 21560 25900 21588 25928
rect 15795 25860 16804 25888
rect 16853 25891 16911 25897
rect 15795 25857 15807 25860
rect 15749 25851 15807 25857
rect 16853 25857 16865 25891
rect 16899 25857 16911 25891
rect 16853 25851 16911 25857
rect 17120 25891 17178 25897
rect 17120 25857 17132 25891
rect 17166 25888 17178 25891
rect 17402 25888 17408 25900
rect 17166 25860 17408 25888
rect 17166 25857 17178 25860
rect 17120 25851 17178 25857
rect 17402 25848 17408 25860
rect 17460 25848 17466 25900
rect 20993 25891 21051 25897
rect 20993 25857 21005 25891
rect 21039 25857 21051 25891
rect 20993 25851 21051 25857
rect 12526 25780 12532 25832
rect 12584 25820 12590 25832
rect 12989 25823 13047 25829
rect 12989 25820 13001 25823
rect 12584 25792 13001 25820
rect 12584 25780 12590 25792
rect 12989 25789 13001 25792
rect 13035 25820 13047 25823
rect 13170 25820 13176 25832
rect 13035 25792 13176 25820
rect 13035 25789 13047 25792
rect 12989 25783 13047 25789
rect 13170 25780 13176 25792
rect 13228 25780 13234 25832
rect 13354 25820 13360 25832
rect 13315 25792 13360 25820
rect 13354 25780 13360 25792
rect 13412 25780 13418 25832
rect 13998 25780 14004 25832
rect 14056 25820 14062 25832
rect 14182 25820 14188 25832
rect 14056 25792 14188 25820
rect 14056 25780 14062 25792
rect 14182 25780 14188 25792
rect 14240 25780 14246 25832
rect 21008 25820 21036 25851
rect 21542 25848 21548 25900
rect 21600 25888 21606 25900
rect 22649 25891 22707 25897
rect 22649 25888 22661 25891
rect 21600 25860 22661 25888
rect 21600 25848 21606 25860
rect 22649 25857 22661 25860
rect 22695 25857 22707 25891
rect 22649 25851 22707 25857
rect 25133 25891 25191 25897
rect 25133 25857 25145 25891
rect 25179 25857 25191 25891
rect 25133 25851 25191 25857
rect 25317 25891 25375 25897
rect 25317 25857 25329 25891
rect 25363 25888 25375 25891
rect 25682 25888 25688 25900
rect 25363 25860 25688 25888
rect 25363 25857 25375 25860
rect 25317 25851 25375 25857
rect 21634 25820 21640 25832
rect 21008 25792 21640 25820
rect 21634 25780 21640 25792
rect 21692 25780 21698 25832
rect 25148 25820 25176 25851
rect 25682 25848 25688 25860
rect 25740 25848 25746 25900
rect 25792 25897 25820 25996
rect 26234 25984 26240 25996
rect 26292 26024 26298 26036
rect 26292 25996 28764 26024
rect 26292 25984 26298 25996
rect 26418 25956 26424 25968
rect 25884 25928 26424 25956
rect 25884 25897 25912 25928
rect 26418 25916 26424 25928
rect 26476 25916 26482 25968
rect 27614 25956 27620 25968
rect 26988 25928 27620 25956
rect 25777 25891 25835 25897
rect 25777 25857 25789 25891
rect 25823 25857 25835 25891
rect 25777 25851 25835 25857
rect 25870 25891 25928 25897
rect 25870 25857 25882 25891
rect 25916 25857 25928 25891
rect 26050 25888 26056 25900
rect 26011 25860 26056 25888
rect 25870 25851 25928 25857
rect 26050 25848 26056 25860
rect 26108 25848 26114 25900
rect 26145 25891 26203 25897
rect 26145 25857 26157 25891
rect 26191 25857 26203 25891
rect 26145 25851 26203 25857
rect 26283 25891 26341 25897
rect 26283 25857 26295 25891
rect 26329 25888 26341 25891
rect 26878 25888 26884 25900
rect 26329 25860 26884 25888
rect 26329 25857 26341 25860
rect 26283 25851 26341 25857
rect 25958 25820 25964 25832
rect 25148 25792 25964 25820
rect 25958 25780 25964 25792
rect 26016 25780 26022 25832
rect 6733 25755 6791 25761
rect 6733 25721 6745 25755
rect 6779 25721 6791 25755
rect 8386 25752 8392 25764
rect 6733 25715 6791 25721
rect 7944 25724 8392 25752
rect 6546 25684 6552 25696
rect 6507 25656 6552 25684
rect 6546 25644 6552 25656
rect 6604 25644 6610 25696
rect 7944 25693 7972 25724
rect 8386 25712 8392 25724
rect 8444 25712 8450 25764
rect 24578 25712 24584 25764
rect 24636 25752 24642 25764
rect 26160 25752 26188 25851
rect 26878 25848 26884 25860
rect 26936 25848 26942 25900
rect 26418 25780 26424 25832
rect 26476 25820 26482 25832
rect 26988 25829 27016 25928
rect 27614 25916 27620 25928
rect 27672 25916 27678 25968
rect 27062 25848 27068 25900
rect 27120 25888 27126 25900
rect 27229 25891 27287 25897
rect 27229 25888 27241 25891
rect 27120 25860 27241 25888
rect 27120 25848 27126 25860
rect 27229 25857 27241 25860
rect 27275 25857 27287 25891
rect 28736 25888 28764 25996
rect 28994 25916 29000 25968
rect 29052 25956 29058 25968
rect 30466 25956 30472 25968
rect 29052 25928 30236 25956
rect 30427 25928 30472 25956
rect 29052 25916 29058 25928
rect 30208 25897 30236 25928
rect 30466 25916 30472 25928
rect 30524 25916 30530 25968
rect 30101 25891 30159 25897
rect 30101 25888 30113 25891
rect 28736 25860 30113 25888
rect 27229 25851 27287 25857
rect 30101 25857 30113 25860
rect 30147 25857 30159 25891
rect 30101 25851 30159 25857
rect 30194 25891 30252 25897
rect 30194 25857 30206 25891
rect 30240 25857 30252 25891
rect 30194 25851 30252 25857
rect 30377 25891 30435 25897
rect 30377 25857 30389 25891
rect 30423 25857 30435 25891
rect 30377 25851 30435 25857
rect 30607 25891 30665 25897
rect 30607 25857 30619 25891
rect 30653 25888 30665 25891
rect 30926 25888 30932 25900
rect 30653 25860 30932 25888
rect 30653 25857 30665 25860
rect 30607 25851 30665 25857
rect 26973 25823 27031 25829
rect 26973 25820 26985 25823
rect 26476 25792 26985 25820
rect 26476 25780 26482 25792
rect 26973 25789 26985 25792
rect 27019 25789 27031 25823
rect 26973 25783 27031 25789
rect 26786 25752 26792 25764
rect 24636 25724 26188 25752
rect 26257 25724 26792 25752
rect 24636 25712 24642 25724
rect 7929 25687 7987 25693
rect 7929 25653 7941 25687
rect 7975 25653 7987 25687
rect 10318 25684 10324 25696
rect 10279 25656 10324 25684
rect 7929 25647 7987 25653
rect 10318 25644 10324 25656
rect 10376 25644 10382 25696
rect 12802 25644 12808 25696
rect 12860 25684 12866 25696
rect 17862 25684 17868 25696
rect 12860 25656 17868 25684
rect 12860 25644 12866 25656
rect 17862 25644 17868 25656
rect 17920 25644 17926 25696
rect 18782 25644 18788 25696
rect 18840 25684 18846 25696
rect 20254 25684 20260 25696
rect 18840 25656 20260 25684
rect 18840 25644 18846 25656
rect 20254 25644 20260 25656
rect 20312 25684 20318 25696
rect 20349 25687 20407 25693
rect 20349 25684 20361 25687
rect 20312 25656 20361 25684
rect 20312 25644 20318 25656
rect 20349 25653 20361 25656
rect 20395 25653 20407 25687
rect 20349 25647 20407 25653
rect 22741 25687 22799 25693
rect 22741 25653 22753 25687
rect 22787 25684 22799 25687
rect 26257 25684 26285 25724
rect 26786 25712 26792 25724
rect 26844 25712 26850 25764
rect 30116 25752 30144 25851
rect 30392 25820 30420 25851
rect 30926 25848 30932 25860
rect 30984 25848 30990 25900
rect 30392 25792 30696 25820
rect 30668 25764 30696 25792
rect 30374 25752 30380 25764
rect 30116 25724 30380 25752
rect 30374 25712 30380 25724
rect 30432 25712 30438 25764
rect 30650 25712 30656 25764
rect 30708 25712 30714 25764
rect 22787 25656 26285 25684
rect 22787 25653 22799 25656
rect 22741 25647 22799 25653
rect 26326 25644 26332 25696
rect 26384 25684 26390 25696
rect 26421 25687 26479 25693
rect 26421 25684 26433 25687
rect 26384 25656 26433 25684
rect 26384 25644 26390 25656
rect 26421 25653 26433 25656
rect 26467 25653 26479 25687
rect 26421 25647 26479 25653
rect 28166 25644 28172 25696
rect 28224 25684 28230 25696
rect 28353 25687 28411 25693
rect 28353 25684 28365 25687
rect 28224 25656 28365 25684
rect 28224 25644 28230 25656
rect 28353 25653 28365 25656
rect 28399 25653 28411 25687
rect 28353 25647 28411 25653
rect 30745 25687 30803 25693
rect 30745 25653 30757 25687
rect 30791 25684 30803 25687
rect 31018 25684 31024 25696
rect 30791 25656 31024 25684
rect 30791 25653 30803 25656
rect 30745 25647 30803 25653
rect 31018 25644 31024 25656
rect 31076 25644 31082 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 5442 25480 5448 25492
rect 5403 25452 5448 25480
rect 5442 25440 5448 25452
rect 5500 25440 5506 25492
rect 9125 25483 9183 25489
rect 9125 25449 9137 25483
rect 9171 25480 9183 25483
rect 9858 25480 9864 25492
rect 9171 25452 9864 25480
rect 9171 25449 9183 25452
rect 9125 25443 9183 25449
rect 9858 25440 9864 25452
rect 9916 25440 9922 25492
rect 10042 25480 10048 25492
rect 10003 25452 10048 25480
rect 10042 25440 10048 25452
rect 10100 25440 10106 25492
rect 10226 25480 10232 25492
rect 10187 25452 10232 25480
rect 10226 25440 10232 25452
rect 10284 25440 10290 25492
rect 10318 25440 10324 25492
rect 10376 25480 10382 25492
rect 10873 25483 10931 25489
rect 10873 25480 10885 25483
rect 10376 25452 10885 25480
rect 10376 25440 10382 25452
rect 10873 25449 10885 25452
rect 10919 25449 10931 25483
rect 10873 25443 10931 25449
rect 11977 25483 12035 25489
rect 11977 25449 11989 25483
rect 12023 25480 12035 25483
rect 12894 25480 12900 25492
rect 12023 25452 12900 25480
rect 12023 25449 12035 25452
rect 11977 25443 12035 25449
rect 12894 25440 12900 25452
rect 12952 25440 12958 25492
rect 17402 25480 17408 25492
rect 17363 25452 17408 25480
rect 17402 25440 17408 25452
rect 17460 25440 17466 25492
rect 18414 25480 18420 25492
rect 17604 25452 18420 25480
rect 14918 25304 14924 25356
rect 14976 25344 14982 25356
rect 15197 25347 15255 25353
rect 15197 25344 15209 25347
rect 14976 25316 15209 25344
rect 14976 25304 14982 25316
rect 15197 25313 15209 25316
rect 15243 25313 15255 25347
rect 15197 25307 15255 25313
rect 5629 25279 5687 25285
rect 5629 25245 5641 25279
rect 5675 25276 5687 25279
rect 6730 25276 6736 25288
rect 5675 25248 6736 25276
rect 5675 25245 5687 25248
rect 5629 25239 5687 25245
rect 6730 25236 6736 25248
rect 6788 25236 6794 25288
rect 6917 25279 6975 25285
rect 6917 25245 6929 25279
rect 6963 25276 6975 25279
rect 8386 25276 8392 25288
rect 6963 25248 8392 25276
rect 6963 25245 6975 25248
rect 6917 25239 6975 25245
rect 8386 25236 8392 25248
rect 8444 25236 8450 25288
rect 8941 25279 8999 25285
rect 8941 25245 8953 25279
rect 8987 25276 8999 25279
rect 9030 25276 9036 25288
rect 8987 25248 9036 25276
rect 8987 25245 8999 25248
rect 8941 25239 8999 25245
rect 9030 25236 9036 25248
rect 9088 25236 9094 25288
rect 11974 25236 11980 25288
rect 12032 25236 12038 25288
rect 12802 25276 12808 25288
rect 12763 25248 12808 25276
rect 12802 25236 12808 25248
rect 12860 25236 12866 25288
rect 15473 25279 15531 25285
rect 15473 25245 15485 25279
rect 15519 25245 15531 25279
rect 15473 25239 15531 25245
rect 16761 25279 16819 25285
rect 16761 25245 16773 25279
rect 16807 25276 16819 25279
rect 17034 25276 17040 25288
rect 16807 25248 17040 25276
rect 16807 25245 16819 25248
rect 16761 25239 16819 25245
rect 9861 25211 9919 25217
rect 9861 25177 9873 25211
rect 9907 25208 9919 25211
rect 10689 25211 10747 25217
rect 10689 25208 10701 25211
rect 9907 25180 10701 25208
rect 9907 25177 9919 25180
rect 9861 25171 9919 25177
rect 10689 25177 10701 25180
rect 10735 25208 10747 25211
rect 10778 25208 10784 25220
rect 10735 25180 10784 25208
rect 10735 25177 10747 25180
rect 10689 25171 10747 25177
rect 10778 25168 10784 25180
rect 10836 25168 10842 25220
rect 11793 25211 11851 25217
rect 11793 25177 11805 25211
rect 11839 25208 11851 25211
rect 11992 25208 12020 25236
rect 15488 25208 15516 25239
rect 17034 25236 17040 25248
rect 17092 25236 17098 25288
rect 17604 25273 17632 25452
rect 18414 25440 18420 25452
rect 18472 25440 18478 25492
rect 19334 25440 19340 25492
rect 19392 25480 19398 25492
rect 21361 25483 21419 25489
rect 19392 25452 20208 25480
rect 19392 25440 19398 25452
rect 17788 25384 18736 25412
rect 17788 25285 17816 25384
rect 17954 25304 17960 25356
rect 18012 25304 18018 25356
rect 17681 25279 17739 25285
rect 17681 25273 17693 25279
rect 17604 25245 17693 25273
rect 17727 25245 17739 25279
rect 17681 25239 17739 25245
rect 17773 25279 17831 25285
rect 17773 25245 17785 25279
rect 17819 25245 17831 25279
rect 17773 25239 17831 25245
rect 17870 25276 17928 25282
rect 17972 25276 18000 25304
rect 17870 25242 17882 25276
rect 17916 25248 18000 25276
rect 18049 25279 18107 25285
rect 17916 25242 17928 25248
rect 17870 25236 17928 25242
rect 18049 25245 18061 25279
rect 18095 25245 18107 25279
rect 18708 25276 18736 25384
rect 19702 25304 19708 25356
rect 19760 25344 19766 25356
rect 19760 25316 19912 25344
rect 19760 25304 19766 25316
rect 19884 25285 19912 25316
rect 19869 25279 19927 25285
rect 18708 25248 19840 25276
rect 18049 25239 18107 25245
rect 16577 25211 16635 25217
rect 16577 25208 16589 25211
rect 11839 25180 12434 25208
rect 15488 25180 16589 25208
rect 11839 25177 11851 25180
rect 11793 25171 11851 25177
rect 6638 25100 6644 25152
rect 6696 25140 6702 25152
rect 6733 25143 6791 25149
rect 6733 25140 6745 25143
rect 6696 25112 6745 25140
rect 6696 25100 6702 25112
rect 6733 25109 6745 25112
rect 6779 25109 6791 25143
rect 6733 25103 6791 25109
rect 9766 25100 9772 25152
rect 9824 25140 9830 25152
rect 10061 25143 10119 25149
rect 10061 25140 10073 25143
rect 9824 25112 10073 25140
rect 9824 25100 9830 25112
rect 10061 25109 10073 25112
rect 10107 25140 10119 25143
rect 10889 25143 10947 25149
rect 10889 25140 10901 25143
rect 10107 25112 10901 25140
rect 10107 25109 10119 25112
rect 10061 25103 10119 25109
rect 10889 25109 10901 25112
rect 10935 25109 10947 25143
rect 11054 25140 11060 25152
rect 11015 25112 11060 25140
rect 10889 25103 10947 25109
rect 11054 25100 11060 25112
rect 11112 25100 11118 25152
rect 11698 25100 11704 25152
rect 11756 25140 11762 25152
rect 11993 25143 12051 25149
rect 11993 25140 12005 25143
rect 11756 25112 12005 25140
rect 11756 25100 11762 25112
rect 11993 25109 12005 25112
rect 12039 25109 12051 25143
rect 12158 25140 12164 25152
rect 12119 25112 12164 25140
rect 11993 25103 12051 25109
rect 12158 25100 12164 25112
rect 12216 25100 12222 25152
rect 12406 25140 12434 25180
rect 16577 25177 16589 25180
rect 16623 25208 16635 25211
rect 16666 25208 16672 25220
rect 16623 25180 16672 25208
rect 16623 25177 16635 25180
rect 16577 25171 16635 25177
rect 16666 25168 16672 25180
rect 16724 25168 16730 25220
rect 18064 25208 18092 25239
rect 18782 25208 18788 25220
rect 18064 25180 18788 25208
rect 18782 25168 18788 25180
rect 18840 25168 18846 25220
rect 19613 25211 19671 25217
rect 19613 25177 19625 25211
rect 19659 25208 19671 25211
rect 19702 25208 19708 25220
rect 19659 25180 19708 25208
rect 19659 25177 19671 25180
rect 19613 25171 19671 25177
rect 19702 25168 19708 25180
rect 19760 25168 19766 25220
rect 19812 25208 19840 25248
rect 19869 25245 19881 25279
rect 19915 25245 19927 25279
rect 19869 25239 19927 25245
rect 19981 25279 20039 25285
rect 19981 25245 19993 25279
rect 20027 25245 20039 25279
rect 19981 25239 20039 25245
rect 20094 25279 20152 25285
rect 20094 25245 20106 25279
rect 20140 25276 20152 25279
rect 20180 25276 20208 25452
rect 21361 25449 21373 25483
rect 21407 25480 21419 25483
rect 22002 25480 22008 25492
rect 21407 25452 22008 25480
rect 21407 25449 21419 25452
rect 21361 25443 21419 25449
rect 22002 25440 22008 25452
rect 22060 25440 22066 25492
rect 26237 25483 26295 25489
rect 26237 25449 26249 25483
rect 26283 25480 26295 25483
rect 27062 25480 27068 25492
rect 26283 25452 27068 25480
rect 26283 25449 26295 25452
rect 26237 25443 26295 25449
rect 27062 25440 27068 25452
rect 27120 25440 27126 25492
rect 26786 25372 26792 25424
rect 26844 25412 26850 25424
rect 30190 25412 30196 25424
rect 26844 25384 30196 25412
rect 26844 25372 26850 25384
rect 30190 25372 30196 25384
rect 30248 25372 30254 25424
rect 25958 25304 25964 25356
rect 26016 25344 26022 25356
rect 31386 25344 31392 25356
rect 26016 25316 28120 25344
rect 26016 25304 26022 25316
rect 20140 25248 20208 25276
rect 20140 25245 20152 25248
rect 20094 25239 20152 25245
rect 19996 25208 20024 25239
rect 20254 25236 20260 25288
rect 20312 25276 20318 25288
rect 21177 25279 21235 25285
rect 20312 25248 20357 25276
rect 20312 25236 20318 25248
rect 21177 25245 21189 25279
rect 21223 25276 21235 25279
rect 21542 25276 21548 25288
rect 21223 25248 21548 25276
rect 21223 25245 21235 25248
rect 21177 25239 21235 25245
rect 21542 25236 21548 25248
rect 21600 25236 21606 25288
rect 22462 25276 22468 25288
rect 22423 25248 22468 25276
rect 22462 25236 22468 25248
rect 22520 25236 22526 25288
rect 22738 25285 22744 25288
rect 22732 25276 22744 25285
rect 22699 25248 22744 25276
rect 22732 25239 22744 25248
rect 22738 25236 22744 25239
rect 22796 25236 22802 25288
rect 24397 25279 24455 25285
rect 24397 25245 24409 25279
rect 24443 25276 24455 25279
rect 26418 25276 26424 25288
rect 24443 25248 26424 25276
rect 24443 25245 24455 25248
rect 24397 25239 24455 25245
rect 26418 25236 26424 25248
rect 26476 25236 26482 25288
rect 26528 25285 26556 25316
rect 26513 25279 26571 25285
rect 26513 25245 26525 25279
rect 26559 25245 26571 25279
rect 26513 25239 26571 25245
rect 26602 25273 26660 25279
rect 26602 25239 26614 25273
rect 26648 25239 26660 25273
rect 26602 25233 26660 25239
rect 26694 25236 26700 25288
rect 26752 25276 26758 25288
rect 26881 25279 26939 25285
rect 26752 25248 26797 25276
rect 26752 25236 26758 25248
rect 26881 25245 26893 25279
rect 26927 25245 26939 25279
rect 26881 25239 26939 25245
rect 19812 25180 20024 25208
rect 12897 25143 12955 25149
rect 12897 25140 12909 25143
rect 12406 25112 12909 25140
rect 12897 25109 12909 25112
rect 12943 25109 12955 25143
rect 12897 25103 12955 25109
rect 16945 25143 17003 25149
rect 16945 25109 16957 25143
rect 16991 25140 17003 25143
rect 17954 25140 17960 25152
rect 16991 25112 17960 25140
rect 16991 25109 17003 25112
rect 16945 25103 17003 25109
rect 17954 25100 17960 25112
rect 18012 25100 18018 25152
rect 19996 25140 20024 25180
rect 24026 25168 24032 25220
rect 24084 25208 24090 25220
rect 24642 25211 24700 25217
rect 24642 25208 24654 25211
rect 24084 25180 24654 25208
rect 24084 25168 24090 25180
rect 24642 25177 24654 25180
rect 24688 25177 24700 25211
rect 24642 25171 24700 25177
rect 24854 25168 24860 25220
rect 24912 25208 24918 25220
rect 24912 25180 26372 25208
rect 24912 25168 24918 25180
rect 20622 25140 20628 25152
rect 19996 25112 20628 25140
rect 20622 25100 20628 25112
rect 20680 25100 20686 25152
rect 23845 25143 23903 25149
rect 23845 25109 23857 25143
rect 23891 25140 23903 25143
rect 24210 25140 24216 25152
rect 23891 25112 24216 25140
rect 23891 25109 23903 25112
rect 23845 25103 23903 25109
rect 24210 25100 24216 25112
rect 24268 25140 24274 25152
rect 24762 25140 24768 25152
rect 24268 25112 24768 25140
rect 24268 25100 24274 25112
rect 24762 25100 24768 25112
rect 24820 25100 24826 25152
rect 25774 25140 25780 25152
rect 25735 25112 25780 25140
rect 25774 25100 25780 25112
rect 25832 25100 25838 25152
rect 26344 25140 26372 25180
rect 26620 25140 26648 25233
rect 26786 25168 26792 25220
rect 26844 25208 26850 25220
rect 26896 25208 26924 25239
rect 27706 25236 27712 25288
rect 27764 25276 27770 25288
rect 27801 25279 27859 25285
rect 27801 25276 27813 25279
rect 27764 25248 27813 25276
rect 27764 25236 27770 25248
rect 27801 25245 27813 25248
rect 27847 25245 27859 25279
rect 27801 25239 27859 25245
rect 27890 25236 27896 25288
rect 27948 25276 27954 25288
rect 28092 25276 28120 25316
rect 30576 25316 31392 25344
rect 28166 25276 28172 25288
rect 27948 25248 27993 25276
rect 28079 25248 28172 25276
rect 27948 25236 27954 25248
rect 28166 25236 28172 25248
rect 28224 25236 28230 25288
rect 28307 25279 28365 25285
rect 28307 25245 28319 25279
rect 28353 25276 28365 25279
rect 29178 25276 29184 25288
rect 28353 25248 29184 25276
rect 28353 25245 28365 25248
rect 28307 25239 28365 25245
rect 29178 25236 29184 25248
rect 29236 25236 29242 25288
rect 30374 25276 30380 25288
rect 30335 25248 30380 25276
rect 30374 25236 30380 25248
rect 30432 25236 30438 25288
rect 30576 25285 30604 25316
rect 31386 25304 31392 25316
rect 31444 25304 31450 25356
rect 30525 25279 30604 25285
rect 30525 25245 30537 25279
rect 30571 25248 30604 25279
rect 30742 25276 30748 25288
rect 30703 25248 30748 25276
rect 30571 25245 30583 25248
rect 30525 25239 30583 25245
rect 30742 25236 30748 25248
rect 30800 25236 30806 25288
rect 30842 25279 30900 25285
rect 30842 25245 30854 25279
rect 30888 25245 30900 25279
rect 30842 25239 30900 25245
rect 26844 25180 26924 25208
rect 28077 25211 28135 25217
rect 26844 25168 26850 25180
rect 28077 25177 28089 25211
rect 28123 25177 28135 25211
rect 30650 25208 30656 25220
rect 30611 25180 30656 25208
rect 28077 25171 28135 25177
rect 26344 25112 26648 25140
rect 26970 25100 26976 25152
rect 27028 25140 27034 25152
rect 28092 25140 28120 25171
rect 30650 25168 30656 25180
rect 30708 25168 30714 25220
rect 27028 25112 28120 25140
rect 28445 25143 28503 25149
rect 27028 25100 27034 25112
rect 28445 25109 28457 25143
rect 28491 25140 28503 25143
rect 28626 25140 28632 25152
rect 28491 25112 28632 25140
rect 28491 25109 28503 25112
rect 28445 25103 28503 25109
rect 28626 25100 28632 25112
rect 28684 25100 28690 25152
rect 28902 25100 28908 25152
rect 28960 25140 28966 25152
rect 30852 25140 30880 25239
rect 28960 25112 30880 25140
rect 31021 25143 31079 25149
rect 28960 25100 28966 25112
rect 31021 25109 31033 25143
rect 31067 25140 31079 25143
rect 33870 25140 33876 25152
rect 31067 25112 33876 25140
rect 31067 25109 31079 25112
rect 31021 25103 31079 25109
rect 33870 25100 33876 25112
rect 33928 25100 33934 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 9582 24936 9588 24948
rect 9543 24908 9588 24936
rect 9582 24896 9588 24908
rect 9640 24896 9646 24948
rect 12894 24936 12900 24948
rect 12855 24908 12900 24936
rect 12894 24896 12900 24908
rect 12952 24896 12958 24948
rect 19058 24936 19064 24948
rect 18892 24908 19064 24936
rect 6914 24868 6920 24880
rect 6875 24840 6920 24868
rect 6914 24828 6920 24840
rect 6972 24828 6978 24880
rect 7117 24871 7175 24877
rect 7117 24868 7129 24871
rect 7116 24837 7129 24868
rect 7163 24837 7175 24871
rect 11054 24868 11060 24880
rect 7116 24831 7175 24837
rect 10888 24840 11060 24868
rect 4706 24800 4712 24812
rect 4667 24772 4712 24800
rect 4706 24760 4712 24772
rect 4764 24760 4770 24812
rect 6178 24760 6184 24812
rect 6236 24800 6242 24812
rect 7116 24800 7144 24831
rect 6236 24772 7144 24800
rect 9769 24803 9827 24809
rect 6236 24760 6242 24772
rect 9769 24769 9781 24803
rect 9815 24800 9827 24803
rect 10888 24800 10916 24840
rect 11054 24828 11060 24840
rect 11112 24828 11118 24880
rect 12158 24868 12164 24880
rect 11164 24840 12164 24868
rect 9815 24772 10916 24800
rect 10965 24803 11023 24809
rect 9815 24769 9827 24772
rect 9769 24763 9827 24769
rect 10965 24769 10977 24803
rect 11011 24800 11023 24803
rect 11164 24800 11192 24840
rect 12158 24828 12164 24840
rect 12216 24828 12222 24880
rect 13538 24828 13544 24880
rect 13596 24868 13602 24880
rect 13596 24840 14044 24868
rect 13596 24828 13602 24840
rect 11773 24803 11831 24809
rect 11773 24800 11785 24803
rect 11011 24772 11192 24800
rect 11256 24772 11785 24800
rect 11011 24769 11023 24772
rect 10965 24763 11023 24769
rect 11256 24732 11284 24772
rect 11773 24769 11785 24772
rect 11819 24769 11831 24803
rect 13630 24800 13636 24812
rect 13591 24772 13636 24800
rect 11773 24763 11831 24769
rect 13630 24760 13636 24772
rect 13688 24760 13694 24812
rect 13725 24803 13783 24809
rect 13725 24769 13737 24803
rect 13771 24769 13783 24803
rect 13725 24763 13783 24769
rect 10796 24704 11284 24732
rect 11517 24735 11575 24741
rect 10796 24673 10824 24704
rect 11517 24701 11529 24735
rect 11563 24701 11575 24735
rect 11517 24695 11575 24701
rect 10781 24667 10839 24673
rect 10781 24633 10793 24667
rect 10827 24633 10839 24667
rect 10781 24627 10839 24633
rect 4525 24599 4583 24605
rect 4525 24565 4537 24599
rect 4571 24596 4583 24599
rect 4614 24596 4620 24608
rect 4571 24568 4620 24596
rect 4571 24565 4583 24568
rect 4525 24559 4583 24565
rect 4614 24556 4620 24568
rect 4672 24556 4678 24608
rect 7098 24596 7104 24608
rect 7059 24568 7104 24596
rect 7098 24556 7104 24568
rect 7156 24556 7162 24608
rect 7282 24596 7288 24608
rect 7243 24568 7288 24596
rect 7282 24556 7288 24568
rect 7340 24556 7346 24608
rect 11532 24596 11560 24695
rect 13354 24692 13360 24744
rect 13412 24732 13418 24744
rect 13740 24732 13768 24763
rect 13814 24760 13820 24812
rect 13872 24800 13878 24812
rect 14016 24809 14044 24840
rect 16666 24828 16672 24880
rect 16724 24868 16730 24880
rect 17865 24871 17923 24877
rect 17865 24868 17877 24871
rect 16724 24840 17877 24868
rect 16724 24828 16730 24840
rect 17865 24837 17877 24840
rect 17911 24868 17923 24871
rect 17911 24840 18184 24868
rect 17911 24837 17923 24840
rect 17865 24831 17923 24837
rect 14001 24803 14059 24809
rect 13872 24772 13917 24800
rect 13872 24760 13878 24772
rect 14001 24769 14013 24803
rect 14047 24800 14059 24803
rect 14274 24800 14280 24812
rect 14047 24772 14280 24800
rect 14047 24769 14059 24772
rect 14001 24763 14059 24769
rect 14274 24760 14280 24772
rect 14332 24760 14338 24812
rect 14912 24803 14970 24809
rect 14912 24769 14924 24803
rect 14958 24800 14970 24803
rect 14958 24772 16712 24800
rect 14958 24769 14970 24772
rect 14912 24763 14970 24769
rect 14458 24732 14464 24744
rect 13412 24704 14464 24732
rect 13412 24692 13418 24704
rect 14458 24692 14464 24704
rect 14516 24692 14522 24744
rect 16684 24741 16712 24772
rect 16850 24760 16856 24812
rect 16908 24800 16914 24812
rect 16945 24803 17003 24809
rect 16945 24800 16957 24803
rect 16908 24772 16957 24800
rect 16908 24760 16914 24772
rect 16945 24769 16957 24772
rect 16991 24769 17003 24803
rect 16945 24763 17003 24769
rect 17037 24803 17095 24809
rect 17037 24769 17049 24803
rect 17083 24769 17095 24803
rect 17037 24763 17095 24769
rect 14645 24735 14703 24741
rect 14645 24701 14657 24735
rect 14691 24701 14703 24735
rect 14645 24695 14703 24701
rect 16669 24735 16727 24741
rect 16669 24701 16681 24735
rect 16715 24701 16727 24735
rect 16669 24695 16727 24701
rect 12836 24636 14136 24664
rect 12836 24596 12864 24636
rect 14108 24608 14136 24636
rect 11532 24568 12864 24596
rect 13357 24599 13415 24605
rect 13357 24565 13369 24599
rect 13403 24596 13415 24599
rect 13998 24596 14004 24608
rect 13403 24568 14004 24596
rect 13403 24565 13415 24568
rect 13357 24559 13415 24565
rect 13998 24556 14004 24568
rect 14056 24556 14062 24608
rect 14090 24556 14096 24608
rect 14148 24596 14154 24608
rect 14660 24596 14688 24695
rect 16758 24692 16764 24744
rect 16816 24732 16822 24744
rect 17052 24732 17080 24763
rect 17126 24760 17132 24812
rect 17184 24800 17190 24812
rect 17313 24803 17371 24809
rect 17184 24772 17229 24800
rect 17184 24760 17190 24772
rect 17313 24769 17325 24803
rect 17359 24800 17371 24803
rect 17770 24800 17776 24812
rect 17359 24772 17776 24800
rect 17359 24769 17371 24772
rect 17313 24763 17371 24769
rect 17770 24760 17776 24772
rect 17828 24760 17834 24812
rect 17954 24760 17960 24812
rect 18012 24800 18018 24812
rect 18049 24803 18107 24809
rect 18049 24800 18061 24803
rect 18012 24772 18061 24800
rect 18012 24760 18018 24772
rect 18049 24769 18061 24772
rect 18095 24769 18107 24803
rect 18156 24800 18184 24840
rect 18892 24809 18920 24908
rect 19058 24896 19064 24908
rect 19116 24936 19122 24948
rect 20714 24936 20720 24948
rect 19116 24908 20720 24936
rect 19116 24896 19122 24908
rect 20714 24896 20720 24908
rect 20772 24896 20778 24948
rect 21085 24939 21143 24945
rect 21085 24905 21097 24939
rect 21131 24936 21143 24939
rect 21174 24936 21180 24948
rect 21131 24908 21180 24936
rect 21131 24905 21143 24908
rect 21085 24899 21143 24905
rect 21174 24896 21180 24908
rect 21232 24896 21238 24948
rect 22094 24896 22100 24948
rect 22152 24936 22158 24948
rect 24026 24936 24032 24948
rect 22152 24908 22784 24936
rect 23987 24908 24032 24936
rect 22152 24896 22158 24908
rect 19978 24877 19984 24880
rect 19972 24868 19984 24877
rect 19352 24840 19840 24868
rect 19939 24840 19984 24868
rect 18693 24803 18751 24809
rect 18693 24800 18705 24803
rect 18156 24772 18705 24800
rect 18049 24763 18107 24769
rect 18693 24769 18705 24772
rect 18739 24769 18751 24803
rect 18693 24763 18751 24769
rect 18877 24803 18935 24809
rect 18877 24769 18889 24803
rect 18923 24769 18935 24803
rect 18877 24763 18935 24769
rect 18966 24760 18972 24812
rect 19024 24800 19030 24812
rect 19352 24800 19380 24840
rect 19024 24772 19380 24800
rect 19024 24760 19030 24772
rect 19426 24760 19432 24812
rect 19484 24800 19490 24812
rect 19705 24803 19763 24809
rect 19705 24800 19717 24803
rect 19484 24772 19717 24800
rect 19484 24760 19490 24772
rect 19705 24769 19717 24772
rect 19751 24769 19763 24803
rect 19812 24800 19840 24840
rect 19972 24831 19984 24840
rect 19978 24828 19984 24831
rect 20036 24828 20042 24880
rect 22554 24868 22560 24880
rect 21836 24840 22560 24868
rect 21836 24800 21864 24840
rect 22554 24828 22560 24840
rect 22612 24828 22618 24880
rect 22756 24877 22784 24908
rect 24026 24896 24032 24908
rect 24084 24896 24090 24948
rect 25774 24936 25780 24948
rect 24320 24908 25780 24936
rect 22741 24871 22799 24877
rect 22741 24837 22753 24871
rect 22787 24837 22799 24871
rect 22741 24831 22799 24837
rect 19812 24772 21864 24800
rect 21913 24803 21971 24809
rect 19705 24763 19763 24769
rect 21913 24769 21925 24803
rect 21959 24800 21971 24803
rect 22646 24800 22652 24812
rect 21959 24772 22652 24800
rect 21959 24769 21971 24772
rect 21913 24763 21971 24769
rect 22646 24760 22652 24772
rect 22704 24760 22710 24812
rect 18233 24735 18291 24741
rect 16816 24704 17448 24732
rect 16816 24692 16822 24704
rect 17310 24664 17316 24676
rect 15580 24636 17316 24664
rect 15580 24596 15608 24636
rect 17310 24624 17316 24636
rect 17368 24624 17374 24676
rect 17420 24664 17448 24704
rect 18233 24701 18245 24735
rect 18279 24732 18291 24735
rect 19334 24732 19340 24744
rect 18279 24704 19340 24732
rect 18279 24701 18291 24704
rect 18233 24695 18291 24701
rect 19334 24692 19340 24704
rect 19392 24692 19398 24744
rect 22756 24732 22784 24831
rect 24320 24809 24348 24908
rect 25774 24896 25780 24908
rect 25832 24896 25838 24948
rect 26329 24939 26387 24945
rect 26329 24905 26341 24939
rect 26375 24936 26387 24939
rect 26694 24936 26700 24948
rect 26375 24908 26700 24936
rect 26375 24905 26387 24908
rect 26329 24899 26387 24905
rect 26694 24896 26700 24908
rect 26752 24896 26758 24948
rect 27890 24896 27896 24948
rect 27948 24936 27954 24948
rect 28353 24939 28411 24945
rect 28353 24936 28365 24939
rect 27948 24908 28365 24936
rect 27948 24896 27954 24908
rect 28353 24905 28365 24908
rect 28399 24905 28411 24939
rect 28353 24899 28411 24905
rect 28997 24939 29055 24945
rect 28997 24905 29009 24939
rect 29043 24936 29055 24939
rect 29178 24936 29184 24948
rect 29043 24908 29184 24936
rect 29043 24905 29055 24908
rect 28997 24899 29055 24905
rect 29178 24896 29184 24908
rect 29236 24896 29242 24948
rect 30466 24896 30472 24948
rect 30524 24896 30530 24948
rect 24854 24868 24860 24880
rect 24412 24840 24860 24868
rect 24412 24809 24440 24840
rect 24854 24828 24860 24840
rect 24912 24828 24918 24880
rect 26602 24828 26608 24880
rect 26660 24868 26666 24880
rect 28902 24868 28908 24880
rect 26660 24840 28908 24868
rect 26660 24828 26666 24840
rect 24305 24803 24363 24809
rect 24305 24769 24317 24803
rect 24351 24769 24363 24803
rect 24305 24763 24363 24769
rect 24397 24803 24455 24809
rect 24397 24769 24409 24803
rect 24443 24769 24455 24803
rect 24397 24763 24455 24769
rect 24486 24760 24492 24812
rect 24544 24800 24550 24812
rect 24670 24800 24676 24812
rect 24544 24772 24589 24800
rect 24631 24772 24676 24800
rect 24544 24760 24550 24772
rect 24670 24760 24676 24772
rect 24728 24760 24734 24812
rect 25225 24803 25283 24809
rect 25225 24769 25237 24803
rect 25271 24769 25283 24803
rect 25958 24800 25964 24812
rect 25919 24772 25964 24800
rect 25225 24763 25283 24769
rect 23014 24732 23020 24744
rect 22756 24704 23020 24732
rect 23014 24692 23020 24704
rect 23072 24732 23078 24744
rect 25240 24732 25268 24763
rect 25958 24760 25964 24772
rect 26016 24760 26022 24812
rect 26145 24803 26203 24809
rect 26145 24769 26157 24803
rect 26191 24800 26203 24803
rect 26786 24800 26792 24812
rect 26191 24772 26792 24800
rect 26191 24769 26203 24772
rect 26145 24763 26203 24769
rect 26786 24760 26792 24772
rect 26844 24760 26850 24812
rect 27062 24760 27068 24812
rect 27120 24800 27126 24812
rect 28828 24809 28856 24840
rect 28902 24828 28908 24840
rect 28960 24828 28966 24880
rect 30190 24828 30196 24880
rect 30248 24868 30254 24880
rect 30484 24868 30512 24896
rect 30248 24840 30788 24868
rect 30248 24828 30254 24840
rect 27229 24803 27287 24809
rect 27229 24800 27241 24803
rect 27120 24772 27241 24800
rect 27120 24760 27126 24772
rect 27229 24769 27241 24772
rect 27275 24769 27287 24803
rect 27229 24763 27287 24769
rect 28813 24803 28871 24809
rect 28813 24769 28825 24803
rect 28859 24769 28871 24803
rect 28813 24763 28871 24769
rect 30377 24803 30435 24809
rect 30377 24769 30389 24803
rect 30423 24769 30435 24803
rect 30377 24763 30435 24769
rect 30469 24803 30527 24809
rect 30469 24769 30481 24803
rect 30515 24769 30527 24803
rect 30469 24763 30527 24769
rect 23072 24704 25268 24732
rect 23072 24692 23078 24704
rect 26418 24692 26424 24744
rect 26476 24732 26482 24744
rect 26973 24735 27031 24741
rect 26973 24732 26985 24735
rect 26476 24704 26985 24732
rect 26476 24692 26482 24704
rect 26973 24701 26985 24704
rect 27019 24701 27031 24735
rect 26973 24695 27031 24701
rect 25130 24664 25136 24676
rect 17420 24636 19656 24664
rect 14148 24568 15608 24596
rect 16025 24599 16083 24605
rect 14148 24556 14154 24568
rect 16025 24565 16037 24599
rect 16071 24596 16083 24599
rect 16850 24596 16856 24608
rect 16071 24568 16856 24596
rect 16071 24565 16083 24568
rect 16025 24559 16083 24565
rect 16850 24556 16856 24568
rect 16908 24556 16914 24608
rect 17954 24556 17960 24608
rect 18012 24596 18018 24608
rect 18966 24596 18972 24608
rect 18012 24568 18972 24596
rect 18012 24556 18018 24568
rect 18966 24556 18972 24568
rect 19024 24556 19030 24608
rect 19061 24599 19119 24605
rect 19061 24565 19073 24599
rect 19107 24596 19119 24599
rect 19518 24596 19524 24608
rect 19107 24568 19524 24596
rect 19107 24565 19119 24568
rect 19061 24559 19119 24565
rect 19518 24556 19524 24568
rect 19576 24556 19582 24608
rect 19628 24596 19656 24636
rect 22112 24636 25136 24664
rect 22112 24605 22140 24636
rect 25130 24624 25136 24636
rect 25188 24624 25194 24676
rect 25409 24667 25467 24673
rect 25409 24633 25421 24667
rect 25455 24664 25467 24667
rect 26510 24664 26516 24676
rect 25455 24636 26516 24664
rect 25455 24633 25467 24636
rect 25409 24627 25467 24633
rect 26510 24624 26516 24636
rect 26568 24664 26574 24676
rect 26878 24664 26884 24676
rect 26568 24636 26884 24664
rect 26568 24624 26574 24636
rect 26878 24624 26884 24636
rect 26936 24624 26942 24676
rect 30392 24664 30420 24763
rect 30484 24732 30512 24763
rect 30558 24760 30564 24812
rect 30616 24800 30622 24812
rect 30760 24809 30788 24840
rect 30745 24803 30803 24809
rect 30616 24772 30661 24800
rect 30616 24760 30622 24772
rect 30745 24769 30757 24803
rect 30791 24769 30803 24803
rect 30745 24763 30803 24769
rect 30834 24760 30840 24812
rect 30892 24800 30898 24812
rect 31205 24803 31263 24809
rect 31205 24800 31217 24803
rect 30892 24772 31217 24800
rect 30892 24760 30898 24772
rect 31205 24769 31217 24772
rect 31251 24769 31263 24803
rect 31386 24800 31392 24812
rect 31205 24763 31263 24769
rect 31312 24772 31392 24800
rect 30650 24732 30656 24744
rect 30484 24704 30656 24732
rect 30650 24692 30656 24704
rect 30708 24692 30714 24744
rect 31312 24732 31340 24772
rect 31386 24760 31392 24772
rect 31444 24760 31450 24812
rect 30760 24704 31340 24732
rect 30760 24664 30788 24704
rect 31202 24664 31208 24676
rect 30392 24636 30788 24664
rect 31163 24636 31208 24664
rect 31202 24624 31208 24636
rect 31260 24624 31266 24676
rect 22097 24599 22155 24605
rect 22097 24596 22109 24599
rect 19628 24568 22109 24596
rect 22097 24565 22109 24568
rect 22143 24565 22155 24599
rect 22097 24559 22155 24565
rect 22738 24556 22744 24608
rect 22796 24596 22802 24608
rect 22833 24599 22891 24605
rect 22833 24596 22845 24599
rect 22796 24568 22845 24596
rect 22796 24556 22802 24568
rect 22833 24565 22845 24568
rect 22879 24565 22891 24599
rect 22833 24559 22891 24565
rect 25958 24556 25964 24608
rect 26016 24596 26022 24608
rect 28994 24596 29000 24608
rect 26016 24568 29000 24596
rect 26016 24556 26022 24568
rect 28994 24556 29000 24568
rect 29052 24556 29058 24608
rect 30101 24599 30159 24605
rect 30101 24565 30113 24599
rect 30147 24596 30159 24599
rect 31110 24596 31116 24608
rect 30147 24568 31116 24596
rect 30147 24565 30159 24568
rect 30101 24559 30159 24565
rect 31110 24556 31116 24568
rect 31168 24556 31174 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 7098 24352 7104 24404
rect 7156 24392 7162 24404
rect 7561 24395 7619 24401
rect 7561 24392 7573 24395
rect 7156 24364 7573 24392
rect 7156 24352 7162 24364
rect 7561 24361 7573 24364
rect 7607 24361 7619 24395
rect 7561 24355 7619 24361
rect 7742 24352 7748 24404
rect 7800 24392 7806 24404
rect 8205 24395 8263 24401
rect 8205 24392 8217 24395
rect 7800 24364 8217 24392
rect 7800 24352 7806 24364
rect 8205 24361 8217 24364
rect 8251 24361 8263 24395
rect 8386 24392 8392 24404
rect 8347 24364 8392 24392
rect 8205 24355 8263 24361
rect 8386 24352 8392 24364
rect 8444 24352 8450 24404
rect 9125 24395 9183 24401
rect 9125 24361 9137 24395
rect 9171 24392 9183 24395
rect 9582 24392 9588 24404
rect 9171 24364 9588 24392
rect 9171 24361 9183 24364
rect 9125 24355 9183 24361
rect 9582 24352 9588 24364
rect 9640 24352 9646 24404
rect 9950 24352 9956 24404
rect 10008 24392 10014 24404
rect 10689 24395 10747 24401
rect 10689 24392 10701 24395
rect 10008 24364 10701 24392
rect 10008 24352 10014 24364
rect 10689 24361 10701 24364
rect 10735 24361 10747 24395
rect 10689 24355 10747 24361
rect 12406 24364 24431 24392
rect 10134 24284 10140 24336
rect 10192 24324 10198 24336
rect 12406 24324 12434 24364
rect 10192 24296 12434 24324
rect 13541 24327 13599 24333
rect 10192 24284 10198 24296
rect 13541 24293 13553 24327
rect 13587 24324 13599 24327
rect 13814 24324 13820 24336
rect 13587 24296 13820 24324
rect 13587 24293 13599 24296
rect 13541 24287 13599 24293
rect 13814 24284 13820 24296
rect 13872 24284 13878 24336
rect 24302 24324 24308 24336
rect 18248 24296 24308 24324
rect 5534 24216 5540 24268
rect 5592 24256 5598 24268
rect 6181 24259 6239 24265
rect 6181 24256 6193 24259
rect 5592 24228 6193 24256
rect 5592 24216 5598 24228
rect 6181 24225 6193 24228
rect 6227 24225 6239 24259
rect 6181 24219 6239 24225
rect 11885 24259 11943 24265
rect 11885 24225 11897 24259
rect 11931 24256 11943 24259
rect 12802 24256 12808 24268
rect 11931 24228 12808 24256
rect 11931 24225 11943 24228
rect 11885 24219 11943 24225
rect 12802 24216 12808 24228
rect 12860 24216 12866 24268
rect 14458 24216 14464 24268
rect 14516 24256 14522 24268
rect 14516 24228 17954 24256
rect 14516 24216 14522 24228
rect 3881 24191 3939 24197
rect 3881 24157 3893 24191
rect 3927 24188 3939 24191
rect 5552 24188 5580 24216
rect 3927 24160 5580 24188
rect 9769 24191 9827 24197
rect 3927 24157 3939 24160
rect 3881 24151 3939 24157
rect 9769 24157 9781 24191
rect 9815 24188 9827 24191
rect 9815 24160 10640 24188
rect 9815 24157 9827 24160
rect 9769 24151 9827 24157
rect 4148 24123 4206 24129
rect 4148 24089 4160 24123
rect 4194 24120 4206 24123
rect 4614 24120 4620 24132
rect 4194 24092 4620 24120
rect 4194 24089 4206 24092
rect 4148 24083 4206 24089
rect 4614 24080 4620 24092
rect 4672 24080 4678 24132
rect 6448 24123 6506 24129
rect 6448 24089 6460 24123
rect 6494 24120 6506 24123
rect 6730 24120 6736 24132
rect 6494 24092 6736 24120
rect 6494 24089 6506 24092
rect 6448 24083 6506 24089
rect 6730 24080 6736 24092
rect 6788 24080 6794 24132
rect 6914 24080 6920 24132
rect 6972 24120 6978 24132
rect 7374 24120 7380 24132
rect 6972 24092 7380 24120
rect 6972 24080 6978 24092
rect 7374 24080 7380 24092
rect 7432 24120 7438 24132
rect 10612 24129 10640 24160
rect 11514 24148 11520 24200
rect 11572 24188 11578 24200
rect 12161 24191 12219 24197
rect 12161 24188 12173 24191
rect 11572 24160 12173 24188
rect 11572 24148 11578 24160
rect 12161 24157 12173 24160
rect 12207 24157 12219 24191
rect 12161 24151 12219 24157
rect 13173 24191 13231 24197
rect 13173 24157 13185 24191
rect 13219 24188 13231 24191
rect 14642 24188 14648 24200
rect 13219 24160 14648 24188
rect 13219 24157 13231 24160
rect 13173 24151 13231 24157
rect 14642 24148 14648 24160
rect 14700 24148 14706 24200
rect 15562 24188 15568 24200
rect 15523 24160 15568 24188
rect 15562 24148 15568 24160
rect 15620 24148 15626 24200
rect 17926 24188 17954 24228
rect 18248 24188 18276 24296
rect 24302 24284 24308 24296
rect 24360 24284 24366 24336
rect 24403 24324 24431 24364
rect 24486 24352 24492 24404
rect 24544 24392 24550 24404
rect 24765 24395 24823 24401
rect 24765 24392 24777 24395
rect 24544 24364 24777 24392
rect 24544 24352 24550 24364
rect 24765 24361 24777 24364
rect 24811 24361 24823 24395
rect 24765 24355 24823 24361
rect 26513 24395 26571 24401
rect 26513 24361 26525 24395
rect 26559 24392 26571 24395
rect 27062 24392 27068 24404
rect 26559 24364 27068 24392
rect 26559 24361 26571 24364
rect 26513 24355 26571 24361
rect 27062 24352 27068 24364
rect 27120 24352 27126 24404
rect 28353 24395 28411 24401
rect 28353 24361 28365 24395
rect 28399 24392 28411 24395
rect 28442 24392 28448 24404
rect 28399 24364 28448 24392
rect 28399 24361 28411 24364
rect 28353 24355 28411 24361
rect 28442 24352 28448 24364
rect 28500 24352 28506 24404
rect 30926 24392 30932 24404
rect 28552 24364 30932 24392
rect 25958 24324 25964 24336
rect 24403 24296 25964 24324
rect 18322 24216 18328 24268
rect 18380 24256 18386 24268
rect 19334 24256 19340 24268
rect 18380 24228 19340 24256
rect 18380 24216 18386 24228
rect 19334 24216 19340 24228
rect 19392 24216 19398 24268
rect 20714 24256 20720 24268
rect 19628 24228 20720 24256
rect 18693 24191 18751 24197
rect 18693 24188 18705 24191
rect 17926 24160 18705 24188
rect 18693 24157 18705 24160
rect 18739 24157 18751 24191
rect 19518 24188 19524 24200
rect 19479 24160 19524 24188
rect 18693 24151 18751 24157
rect 19518 24148 19524 24160
rect 19576 24148 19582 24200
rect 19628 24197 19656 24228
rect 20714 24216 20720 24228
rect 20772 24216 20778 24268
rect 21361 24259 21419 24265
rect 21361 24225 21373 24259
rect 21407 24256 21419 24259
rect 23198 24256 23204 24268
rect 21407 24228 23204 24256
rect 21407 24225 21419 24228
rect 21361 24219 21419 24225
rect 23198 24216 23204 24228
rect 23256 24216 23262 24268
rect 19613 24191 19671 24197
rect 19613 24157 19625 24191
rect 19659 24157 19671 24191
rect 19613 24151 19671 24157
rect 19702 24148 19708 24200
rect 19760 24188 19766 24200
rect 19889 24191 19947 24197
rect 19760 24160 19805 24188
rect 19760 24148 19766 24160
rect 19889 24157 19901 24191
rect 19935 24188 19947 24191
rect 19978 24188 19984 24200
rect 19935 24160 19984 24188
rect 19935 24157 19947 24160
rect 19889 24151 19947 24157
rect 19978 24148 19984 24160
rect 20036 24188 20042 24200
rect 20254 24188 20260 24200
rect 20036 24160 20260 24188
rect 20036 24148 20042 24160
rect 20254 24148 20260 24160
rect 20312 24148 20318 24200
rect 20441 24191 20499 24197
rect 20441 24157 20453 24191
rect 20487 24188 20499 24191
rect 21542 24188 21548 24200
rect 20487 24160 21548 24188
rect 20487 24157 20499 24160
rect 20441 24151 20499 24157
rect 21542 24148 21548 24160
rect 21600 24188 21606 24200
rect 21919 24191 21977 24197
rect 21600 24185 21864 24188
rect 21919 24185 21931 24191
rect 21600 24160 21931 24185
rect 21600 24148 21606 24160
rect 21836 24157 21931 24160
rect 21965 24185 21977 24191
rect 22094 24188 22100 24200
rect 22020 24185 22100 24188
rect 21965 24160 22100 24185
rect 21965 24157 22048 24160
rect 21919 24151 21977 24157
rect 22094 24148 22100 24160
rect 22152 24148 22158 24200
rect 24403 24197 24431 24296
rect 25958 24284 25964 24296
rect 26016 24284 26022 24336
rect 26878 24284 26884 24336
rect 26936 24324 26942 24336
rect 28552 24324 28580 24364
rect 30926 24352 30932 24364
rect 30984 24352 30990 24404
rect 31386 24352 31392 24404
rect 31444 24392 31450 24404
rect 32769 24395 32827 24401
rect 32769 24392 32781 24395
rect 31444 24364 32781 24392
rect 31444 24352 31450 24364
rect 32769 24361 32781 24364
rect 32815 24361 32827 24395
rect 32769 24355 32827 24361
rect 26936 24296 28580 24324
rect 26936 24284 26942 24296
rect 26053 24259 26111 24265
rect 26053 24225 26065 24259
rect 26099 24256 26111 24259
rect 28902 24256 28908 24268
rect 26099 24228 27016 24256
rect 26099 24225 26111 24228
rect 26053 24219 26111 24225
rect 23109 24191 23167 24197
rect 23109 24157 23121 24191
rect 23155 24188 23167 24191
rect 24397 24191 24455 24197
rect 23155 24160 24348 24188
rect 23155 24157 23167 24160
rect 23109 24151 23167 24157
rect 8021 24123 8079 24129
rect 8021 24120 8033 24123
rect 7432 24092 8033 24120
rect 7432 24080 7438 24092
rect 8021 24089 8033 24092
rect 8067 24120 8079 24123
rect 8941 24123 8999 24129
rect 8941 24120 8953 24123
rect 8067 24092 8953 24120
rect 8067 24089 8079 24092
rect 8021 24083 8079 24089
rect 8941 24089 8953 24092
rect 8987 24089 8999 24123
rect 8941 24083 8999 24089
rect 10597 24123 10655 24129
rect 10597 24089 10609 24123
rect 10643 24120 10655 24123
rect 11790 24120 11796 24132
rect 10643 24092 11796 24120
rect 10643 24089 10655 24092
rect 10597 24083 10655 24089
rect 11790 24080 11796 24092
rect 11848 24080 11854 24132
rect 13357 24123 13415 24129
rect 13357 24089 13369 24123
rect 13403 24120 13415 24123
rect 16206 24120 16212 24132
rect 13403 24092 16212 24120
rect 13403 24089 13415 24092
rect 13357 24083 13415 24089
rect 16206 24080 16212 24092
rect 16264 24080 16270 24132
rect 17310 24120 17316 24132
rect 17271 24092 17316 24120
rect 17310 24080 17316 24092
rect 17368 24080 17374 24132
rect 18509 24123 18567 24129
rect 18509 24089 18521 24123
rect 18555 24120 18567 24123
rect 20622 24120 20628 24132
rect 18555 24092 19564 24120
rect 20583 24092 20628 24120
rect 18555 24089 18567 24092
rect 18509 24083 18567 24089
rect 5261 24055 5319 24061
rect 5261 24021 5273 24055
rect 5307 24052 5319 24055
rect 5350 24052 5356 24064
rect 5307 24024 5356 24052
rect 5307 24021 5319 24024
rect 5261 24015 5319 24021
rect 5350 24012 5356 24024
rect 5408 24012 5414 24064
rect 6178 24012 6184 24064
rect 6236 24052 6242 24064
rect 8221 24055 8279 24061
rect 8221 24052 8233 24055
rect 6236 24024 8233 24052
rect 6236 24012 6242 24024
rect 8221 24021 8233 24024
rect 8267 24052 8279 24055
rect 8570 24052 8576 24064
rect 8267 24024 8576 24052
rect 8267 24021 8279 24024
rect 8221 24015 8279 24021
rect 8570 24012 8576 24024
rect 8628 24052 8634 24064
rect 9030 24052 9036 24064
rect 8628 24024 9036 24052
rect 8628 24012 8634 24024
rect 9030 24012 9036 24024
rect 9088 24052 9094 24064
rect 9141 24055 9199 24061
rect 9141 24052 9153 24055
rect 9088 24024 9153 24052
rect 9088 24012 9094 24024
rect 9141 24021 9153 24024
rect 9187 24021 9199 24055
rect 9306 24052 9312 24064
rect 9267 24024 9312 24052
rect 9141 24015 9199 24021
rect 9306 24012 9312 24024
rect 9364 24012 9370 24064
rect 9953 24055 10011 24061
rect 9953 24021 9965 24055
rect 9999 24052 10011 24055
rect 10134 24052 10140 24064
rect 9999 24024 10140 24052
rect 9999 24021 10011 24024
rect 9953 24015 10011 24021
rect 10134 24012 10140 24024
rect 10192 24012 10198 24064
rect 19288 24061 19294 24064
rect 19245 24055 19294 24061
rect 19245 24021 19257 24055
rect 19291 24021 19294 24055
rect 19245 24015 19294 24021
rect 19288 24012 19294 24015
rect 19346 24052 19352 24064
rect 19536 24052 19564 24092
rect 20622 24080 20628 24092
rect 20680 24080 20686 24132
rect 21174 24120 21180 24132
rect 21087 24092 21180 24120
rect 21174 24080 21180 24092
rect 21232 24120 21238 24132
rect 21634 24120 21640 24132
rect 21232 24092 21640 24120
rect 21232 24080 21238 24092
rect 21634 24080 21640 24092
rect 21692 24080 21698 24132
rect 22646 24080 22652 24132
rect 22704 24120 22710 24132
rect 22925 24123 22983 24129
rect 22925 24120 22937 24123
rect 22704 24092 22937 24120
rect 22704 24080 22710 24092
rect 22925 24089 22937 24092
rect 22971 24120 22983 24123
rect 23661 24123 23719 24129
rect 23661 24120 23673 24123
rect 22971 24092 23673 24120
rect 22971 24089 22983 24092
rect 22925 24083 22983 24089
rect 23661 24089 23673 24092
rect 23707 24089 23719 24123
rect 24320 24120 24348 24160
rect 24397 24157 24409 24191
rect 24443 24157 24455 24191
rect 24854 24188 24860 24200
rect 24397 24151 24455 24157
rect 24505 24160 24860 24188
rect 24505 24120 24533 24160
rect 24854 24148 24860 24160
rect 24912 24148 24918 24200
rect 25038 24148 25044 24200
rect 25096 24188 25102 24200
rect 25685 24191 25743 24197
rect 25685 24188 25697 24191
rect 25096 24160 25697 24188
rect 25096 24148 25102 24160
rect 25685 24157 25697 24160
rect 25731 24157 25743 24191
rect 26786 24188 26792 24200
rect 26747 24160 26792 24188
rect 25685 24151 25743 24157
rect 26786 24148 26792 24160
rect 26844 24148 26850 24200
rect 26988 24197 27016 24228
rect 28368 24228 28908 24256
rect 28368 24197 28396 24228
rect 28902 24216 28908 24228
rect 28960 24216 28966 24268
rect 31110 24216 31116 24268
rect 31168 24256 31174 24268
rect 31168 24228 31524 24256
rect 31168 24216 31174 24228
rect 26878 24188 26936 24194
rect 26878 24154 26890 24188
rect 26924 24154 26936 24188
rect 26878 24148 26936 24154
rect 26973 24191 27031 24197
rect 26973 24157 26985 24191
rect 27019 24157 27031 24191
rect 26973 24151 27031 24157
rect 27157 24191 27215 24197
rect 27157 24157 27169 24191
rect 27203 24157 27215 24191
rect 27157 24151 27215 24157
rect 28353 24191 28411 24197
rect 28353 24157 28365 24191
rect 28399 24157 28411 24191
rect 28353 24151 28411 24157
rect 24320 24092 24533 24120
rect 24581 24123 24639 24129
rect 23661 24083 23719 24089
rect 24581 24089 24593 24123
rect 24627 24120 24639 24123
rect 25314 24120 25320 24132
rect 24627 24092 25320 24120
rect 24627 24089 24639 24092
rect 24581 24083 24639 24089
rect 25314 24080 25320 24092
rect 25372 24080 25378 24132
rect 25869 24123 25927 24129
rect 25869 24089 25881 24123
rect 25915 24120 25927 24123
rect 26142 24120 26148 24132
rect 25915 24092 26148 24120
rect 25915 24089 25927 24092
rect 25869 24083 25927 24089
rect 26142 24080 26148 24092
rect 26200 24080 26206 24132
rect 26694 24080 26700 24132
rect 26752 24120 26758 24132
rect 26893 24120 26921 24148
rect 26752 24092 26921 24120
rect 26752 24080 26758 24092
rect 21192 24052 21220 24080
rect 19346 24024 19393 24052
rect 19536 24024 21220 24052
rect 22097 24055 22155 24061
rect 19346 24012 19352 24024
rect 22097 24021 22109 24055
rect 22143 24052 22155 24055
rect 22830 24052 22836 24064
rect 22143 24024 22836 24052
rect 22143 24021 22155 24024
rect 22097 24015 22155 24021
rect 22830 24012 22836 24024
rect 22888 24012 22894 24064
rect 23750 24052 23756 24064
rect 23711 24024 23756 24052
rect 23750 24012 23756 24024
rect 23808 24012 23814 24064
rect 25682 24012 25688 24064
rect 25740 24052 25746 24064
rect 27172 24052 27200 24151
rect 28442 24148 28448 24200
rect 28500 24188 28506 24200
rect 28537 24191 28595 24197
rect 28537 24188 28549 24191
rect 28500 24160 28549 24188
rect 28500 24148 28506 24160
rect 28537 24157 28549 24160
rect 28583 24157 28595 24191
rect 28537 24151 28595 24157
rect 29549 24191 29607 24197
rect 29549 24157 29561 24191
rect 29595 24188 29607 24191
rect 30098 24188 30104 24200
rect 29595 24160 30104 24188
rect 29595 24157 29607 24160
rect 29549 24151 29607 24157
rect 30098 24148 30104 24160
rect 30156 24188 30162 24200
rect 31389 24191 31447 24197
rect 31389 24188 31401 24191
rect 30156 24160 31401 24188
rect 30156 24148 30162 24160
rect 31389 24157 31401 24160
rect 31435 24157 31447 24191
rect 31496 24188 31524 24228
rect 31645 24191 31703 24197
rect 31645 24188 31657 24191
rect 31496 24160 31657 24188
rect 31389 24151 31447 24157
rect 31645 24157 31657 24160
rect 31691 24157 31703 24191
rect 31645 24151 31703 24157
rect 28258 24080 28264 24132
rect 28316 24120 28322 24132
rect 29794 24123 29852 24129
rect 29794 24120 29806 24123
rect 28316 24092 29806 24120
rect 28316 24080 28322 24092
rect 29794 24089 29806 24092
rect 29840 24089 29852 24123
rect 29794 24083 29852 24089
rect 28350 24052 28356 24064
rect 25740 24024 28356 24052
rect 25740 24012 25746 24024
rect 28350 24012 28356 24024
rect 28408 24052 28414 24064
rect 28718 24052 28724 24064
rect 28408 24024 28724 24052
rect 28408 24012 28414 24024
rect 28718 24012 28724 24024
rect 28776 24012 28782 24064
rect 30282 24012 30288 24064
rect 30340 24052 30346 24064
rect 30929 24055 30987 24061
rect 30929 24052 30941 24055
rect 30340 24024 30941 24052
rect 30340 24012 30346 24024
rect 30929 24021 30941 24024
rect 30975 24021 30987 24055
rect 30929 24015 30987 24021
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 4706 23808 4712 23860
rect 4764 23848 4770 23860
rect 5537 23851 5595 23857
rect 5537 23848 5549 23851
rect 4764 23820 5549 23848
rect 4764 23808 4770 23820
rect 5537 23817 5549 23820
rect 5583 23817 5595 23851
rect 6914 23848 6920 23860
rect 5537 23811 5595 23817
rect 6288 23820 6920 23848
rect 5169 23783 5227 23789
rect 5169 23749 5181 23783
rect 5215 23749 5227 23783
rect 5169 23743 5227 23749
rect 5385 23783 5443 23789
rect 5385 23749 5397 23783
rect 5431 23780 5443 23783
rect 6178 23780 6184 23792
rect 5431 23752 6184 23780
rect 5431 23749 5443 23752
rect 5385 23743 5443 23749
rect 4525 23715 4583 23721
rect 4525 23681 4537 23715
rect 4571 23712 4583 23715
rect 4890 23712 4896 23724
rect 4571 23684 4896 23712
rect 4571 23681 4583 23684
rect 4525 23675 4583 23681
rect 4890 23672 4896 23684
rect 4948 23672 4954 23724
rect 5184 23712 5212 23743
rect 6178 23740 6184 23752
rect 6236 23740 6242 23792
rect 6288 23712 6316 23820
rect 6914 23808 6920 23820
rect 6972 23808 6978 23860
rect 7742 23848 7748 23860
rect 7703 23820 7748 23848
rect 7742 23808 7748 23820
rect 7800 23808 7806 23860
rect 9582 23848 9588 23860
rect 9543 23820 9588 23848
rect 9582 23808 9588 23820
rect 9640 23808 9646 23860
rect 10778 23848 10784 23860
rect 10428 23820 10784 23848
rect 10428 23789 10456 23820
rect 10778 23808 10784 23820
rect 10836 23848 10842 23860
rect 11514 23848 11520 23860
rect 10836 23820 11520 23848
rect 10836 23808 10842 23820
rect 11514 23808 11520 23820
rect 11572 23808 11578 23860
rect 12069 23851 12127 23857
rect 12069 23817 12081 23851
rect 12115 23848 12127 23851
rect 17126 23848 17132 23860
rect 12115 23820 17132 23848
rect 12115 23817 12127 23820
rect 12069 23811 12127 23817
rect 17126 23808 17132 23820
rect 17184 23808 17190 23860
rect 17236 23820 22784 23848
rect 10413 23783 10471 23789
rect 6380 23752 8248 23780
rect 6380 23721 6408 23752
rect 6638 23721 6644 23724
rect 5184 23684 6316 23712
rect 6365 23715 6423 23721
rect 6365 23681 6377 23715
rect 6411 23681 6423 23715
rect 6632 23712 6644 23721
rect 6599 23684 6644 23712
rect 6365 23675 6423 23681
rect 6632 23675 6644 23684
rect 6638 23672 6644 23675
rect 6696 23672 6702 23724
rect 8220 23721 8248 23752
rect 10413 23749 10425 23783
rect 10459 23749 10471 23783
rect 10413 23743 10471 23749
rect 10629 23783 10687 23789
rect 10629 23749 10641 23783
rect 10675 23780 10687 23783
rect 11698 23780 11704 23792
rect 10675 23752 11704 23780
rect 10675 23749 10687 23752
rect 10629 23743 10687 23749
rect 11698 23740 11704 23752
rect 11756 23740 11762 23792
rect 13998 23740 14004 23792
rect 14056 23780 14062 23792
rect 14338 23783 14396 23789
rect 14338 23780 14350 23783
rect 14056 23752 14350 23780
rect 14056 23740 14062 23752
rect 14338 23749 14350 23752
rect 14384 23749 14396 23783
rect 14338 23743 14396 23749
rect 14642 23740 14648 23792
rect 14700 23780 14706 23792
rect 16945 23783 17003 23789
rect 16945 23780 16957 23783
rect 14700 23752 16957 23780
rect 14700 23740 14706 23752
rect 16945 23749 16957 23752
rect 16991 23780 17003 23783
rect 17236 23780 17264 23820
rect 16991 23752 17264 23780
rect 16991 23749 17003 23752
rect 16945 23743 17003 23749
rect 17310 23740 17316 23792
rect 17368 23780 17374 23792
rect 19518 23789 19524 23792
rect 19490 23783 19524 23789
rect 17368 23752 19288 23780
rect 17368 23740 17374 23752
rect 13351 23724 13357 23727
rect 8205 23715 8263 23721
rect 8205 23681 8217 23715
rect 8251 23712 8263 23715
rect 8294 23712 8300 23724
rect 8251 23684 8300 23712
rect 8251 23681 8263 23684
rect 8205 23675 8263 23681
rect 8294 23672 8300 23684
rect 8352 23672 8358 23724
rect 8478 23721 8484 23724
rect 8472 23675 8484 23721
rect 8536 23712 8542 23724
rect 8536 23684 8572 23712
rect 8478 23672 8484 23675
rect 8536 23672 8542 23684
rect 11422 23672 11428 23724
rect 11480 23712 11486 23724
rect 11885 23715 11943 23721
rect 11885 23712 11897 23715
rect 11480 23684 11897 23712
rect 11480 23672 11486 23684
rect 11885 23681 11897 23684
rect 11931 23681 11943 23715
rect 11885 23675 11943 23681
rect 13245 23715 13303 23721
rect 13245 23681 13257 23715
rect 13291 23681 13303 23715
rect 13245 23675 13303 23681
rect 13338 23718 13357 23724
rect 13338 23684 13350 23718
rect 13338 23678 13357 23684
rect 13351 23675 13357 23678
rect 13409 23675 13415 23727
rect 13470 23715 13528 23721
rect 13470 23681 13482 23715
rect 13516 23712 13528 23715
rect 13633 23715 13691 23721
rect 13516 23684 13584 23712
rect 13516 23681 13528 23684
rect 13470 23675 13528 23681
rect 13260 23644 13288 23675
rect 13556 23644 13584 23684
rect 13633 23681 13645 23715
rect 13679 23712 13691 23715
rect 13906 23712 13912 23724
rect 13679 23684 13912 23712
rect 13679 23681 13691 23684
rect 13633 23675 13691 23681
rect 13906 23672 13912 23684
rect 13964 23672 13970 23724
rect 14090 23712 14096 23724
rect 14051 23684 14096 23712
rect 14090 23672 14096 23684
rect 14148 23672 14154 23724
rect 17420 23721 17448 23752
rect 16761 23715 16819 23721
rect 16761 23681 16773 23715
rect 16807 23681 16819 23715
rect 16761 23675 16819 23681
rect 17405 23715 17463 23721
rect 17405 23681 17417 23715
rect 17451 23681 17463 23715
rect 17405 23675 17463 23681
rect 13998 23644 14004 23656
rect 13260 23616 13397 23644
rect 13556 23616 14004 23644
rect 13262 23536 13268 23588
rect 13320 23576 13326 23588
rect 13369 23576 13397 23616
rect 13998 23604 14004 23616
rect 14056 23604 14062 23656
rect 13320 23548 13397 23576
rect 15473 23579 15531 23585
rect 13320 23536 13326 23548
rect 15473 23545 15485 23579
rect 15519 23576 15531 23579
rect 16206 23576 16212 23588
rect 15519 23548 16212 23576
rect 15519 23545 15531 23548
rect 15473 23539 15531 23545
rect 16206 23536 16212 23548
rect 16264 23536 16270 23588
rect 4341 23511 4399 23517
rect 4341 23477 4353 23511
rect 4387 23508 4399 23511
rect 4614 23508 4620 23520
rect 4387 23480 4620 23508
rect 4387 23477 4399 23480
rect 4341 23471 4399 23477
rect 4614 23468 4620 23480
rect 4672 23468 4678 23520
rect 5350 23508 5356 23520
rect 5311 23480 5356 23508
rect 5350 23468 5356 23480
rect 5408 23468 5414 23520
rect 10594 23508 10600 23520
rect 10555 23480 10600 23508
rect 10594 23468 10600 23480
rect 10652 23468 10658 23520
rect 10778 23508 10784 23520
rect 10739 23480 10784 23508
rect 10778 23468 10784 23480
rect 10836 23468 10842 23520
rect 12989 23511 13047 23517
rect 12989 23477 13001 23511
rect 13035 23508 13047 23511
rect 13078 23508 13084 23520
rect 13035 23480 13084 23508
rect 13035 23477 13047 23480
rect 12989 23471 13047 23477
rect 13078 23468 13084 23480
rect 13136 23468 13142 23520
rect 16776 23508 16804 23675
rect 17494 23672 17500 23724
rect 17552 23712 17558 23724
rect 19260 23721 19288 23752
rect 19490 23749 19502 23783
rect 19490 23743 19524 23749
rect 19518 23740 19524 23743
rect 19576 23740 19582 23792
rect 19978 23740 19984 23792
rect 20036 23780 20042 23792
rect 22554 23780 22560 23792
rect 20036 23752 22560 23780
rect 20036 23740 20042 23752
rect 22554 23740 22560 23752
rect 22612 23740 22618 23792
rect 22756 23780 22784 23820
rect 22830 23808 22836 23860
rect 22888 23848 22894 23860
rect 23290 23848 23296 23860
rect 22888 23820 23296 23848
rect 22888 23808 22894 23820
rect 23290 23808 23296 23820
rect 23348 23808 23354 23860
rect 25041 23851 25099 23857
rect 25041 23817 25053 23851
rect 25087 23848 25099 23851
rect 25130 23848 25136 23860
rect 25087 23820 25136 23848
rect 25087 23817 25099 23820
rect 25041 23811 25099 23817
rect 25130 23808 25136 23820
rect 25188 23808 25194 23860
rect 25774 23808 25780 23860
rect 25832 23848 25838 23860
rect 26050 23848 26056 23860
rect 25832 23820 26056 23848
rect 25832 23808 25838 23820
rect 26050 23808 26056 23820
rect 26108 23808 26114 23860
rect 28258 23848 28264 23860
rect 28219 23820 28264 23848
rect 28258 23808 28264 23820
rect 28316 23808 28322 23860
rect 28718 23808 28724 23860
rect 28776 23808 28782 23860
rect 29825 23851 29883 23857
rect 29825 23817 29837 23851
rect 29871 23848 29883 23851
rect 30558 23848 30564 23860
rect 29871 23820 30564 23848
rect 29871 23817 29883 23820
rect 29825 23811 29883 23817
rect 30558 23808 30564 23820
rect 30616 23808 30622 23860
rect 22756 23752 24256 23780
rect 17661 23715 17719 23721
rect 17661 23712 17673 23715
rect 17552 23684 17673 23712
rect 17552 23672 17558 23684
rect 17661 23681 17673 23684
rect 17707 23681 17719 23715
rect 17661 23675 17719 23681
rect 19245 23715 19303 23721
rect 19245 23681 19257 23715
rect 19291 23681 19303 23715
rect 22094 23712 22100 23724
rect 22055 23684 22100 23712
rect 19245 23675 19303 23681
rect 22094 23672 22100 23684
rect 22152 23672 22158 23724
rect 22646 23672 22652 23724
rect 22704 23712 22710 23724
rect 23201 23715 23259 23721
rect 23201 23712 23213 23715
rect 22704 23684 23213 23712
rect 22704 23672 22710 23684
rect 23201 23681 23213 23684
rect 23247 23681 23259 23715
rect 24228 23712 24256 23752
rect 24302 23740 24308 23792
rect 24360 23780 24366 23792
rect 26694 23780 26700 23792
rect 24360 23752 26700 23780
rect 24360 23740 24366 23752
rect 25038 23712 25044 23724
rect 24228 23684 25044 23712
rect 23201 23675 23259 23681
rect 25038 23672 25044 23684
rect 25096 23672 25102 23724
rect 25314 23712 25320 23724
rect 25227 23684 25320 23712
rect 25314 23672 25320 23684
rect 25372 23672 25378 23724
rect 25424 23721 25452 23752
rect 26694 23740 26700 23752
rect 26752 23780 26758 23792
rect 28736 23780 28764 23808
rect 26752 23752 28672 23780
rect 28736 23752 28948 23780
rect 26752 23740 26758 23752
rect 25409 23715 25467 23721
rect 25409 23681 25421 23715
rect 25455 23681 25467 23715
rect 25409 23675 25467 23681
rect 25498 23672 25504 23724
rect 25556 23712 25562 23724
rect 25556 23684 25601 23712
rect 25556 23672 25562 23684
rect 25682 23672 25688 23724
rect 25740 23712 25746 23724
rect 26142 23712 26148 23724
rect 25740 23684 25785 23712
rect 26055 23684 26148 23712
rect 25740 23672 25746 23684
rect 26142 23672 26148 23684
rect 26200 23672 26206 23724
rect 26329 23715 26387 23721
rect 26329 23681 26341 23715
rect 26375 23712 26387 23715
rect 26418 23712 26424 23724
rect 26375 23684 26424 23712
rect 26375 23681 26387 23684
rect 26329 23675 26387 23681
rect 26418 23672 26424 23684
rect 26476 23672 26482 23724
rect 27890 23712 27896 23724
rect 26528 23684 27896 23712
rect 20990 23604 20996 23656
rect 21048 23644 21054 23656
rect 21821 23647 21879 23653
rect 21821 23644 21833 23647
rect 21048 23616 21833 23644
rect 21048 23604 21054 23616
rect 21821 23613 21833 23616
rect 21867 23613 21879 23647
rect 25332 23644 25360 23672
rect 25866 23644 25872 23656
rect 25332 23616 25872 23644
rect 21821 23607 21879 23613
rect 25866 23604 25872 23616
rect 25924 23604 25930 23656
rect 26160 23644 26188 23672
rect 26528 23644 26556 23684
rect 27890 23672 27896 23684
rect 27948 23672 27954 23724
rect 28074 23672 28080 23724
rect 28132 23712 28138 23724
rect 28258 23712 28264 23724
rect 28132 23684 28264 23712
rect 28132 23672 28138 23684
rect 28258 23672 28264 23684
rect 28316 23672 28322 23724
rect 28644 23721 28672 23752
rect 28517 23715 28575 23721
rect 28517 23681 28529 23715
rect 28563 23712 28575 23715
rect 28629 23715 28687 23721
rect 28563 23681 28580 23712
rect 28517 23675 28580 23681
rect 28629 23681 28641 23715
rect 28675 23681 28687 23715
rect 28629 23675 28687 23681
rect 26160 23616 26556 23644
rect 28552 23644 28580 23675
rect 28718 23672 28724 23724
rect 28776 23712 28782 23724
rect 28920 23721 28948 23752
rect 30282 23740 30288 23792
rect 30340 23780 30346 23792
rect 30745 23783 30803 23789
rect 30340 23752 30512 23780
rect 30340 23740 30346 23752
rect 28905 23715 28963 23721
rect 28776 23684 28821 23712
rect 28776 23672 28782 23684
rect 28905 23681 28917 23715
rect 28951 23681 28963 23715
rect 28905 23675 28963 23681
rect 28994 23672 29000 23724
rect 29052 23712 29058 23724
rect 29457 23715 29515 23721
rect 29457 23712 29469 23715
rect 29052 23684 29469 23712
rect 29052 23672 29058 23684
rect 29457 23681 29469 23684
rect 29503 23681 29515 23715
rect 29457 23675 29515 23681
rect 29641 23715 29699 23721
rect 29641 23681 29653 23715
rect 29687 23681 29699 23715
rect 29641 23675 29699 23681
rect 29656 23644 29684 23675
rect 29730 23672 29736 23724
rect 29788 23712 29794 23724
rect 30374 23712 30380 23724
rect 29788 23684 30380 23712
rect 29788 23672 29794 23684
rect 30374 23672 30380 23684
rect 30432 23672 30438 23724
rect 30484 23721 30512 23752
rect 30745 23749 30757 23783
rect 30791 23780 30803 23783
rect 31386 23780 31392 23792
rect 30791 23752 31392 23780
rect 30791 23749 30803 23752
rect 30745 23743 30803 23749
rect 31386 23740 31392 23752
rect 31444 23740 31450 23792
rect 30470 23715 30528 23721
rect 30470 23681 30482 23715
rect 30516 23681 30528 23715
rect 30470 23675 30528 23681
rect 28552 23616 30420 23644
rect 30392 23588 30420 23616
rect 18785 23579 18843 23585
rect 18785 23545 18797 23579
rect 18831 23576 18843 23579
rect 18874 23576 18880 23588
rect 18831 23548 18880 23576
rect 18831 23545 18843 23548
rect 18785 23539 18843 23545
rect 18874 23536 18880 23548
rect 18932 23536 18938 23588
rect 20438 23536 20444 23588
rect 20496 23576 20502 23588
rect 20625 23579 20683 23585
rect 20625 23576 20637 23579
rect 20496 23548 20637 23576
rect 20496 23536 20502 23548
rect 20625 23545 20637 23548
rect 20671 23545 20683 23579
rect 20625 23539 20683 23545
rect 22094 23536 22100 23588
rect 22152 23576 22158 23588
rect 22278 23576 22284 23588
rect 22152 23548 22284 23576
rect 22152 23536 22158 23548
rect 22278 23536 22284 23548
rect 22336 23536 22342 23588
rect 24394 23536 24400 23588
rect 24452 23576 24458 23588
rect 26145 23579 26203 23585
rect 26145 23576 26157 23579
rect 24452 23548 26157 23576
rect 24452 23536 24458 23548
rect 26145 23545 26157 23548
rect 26191 23545 26203 23579
rect 26145 23539 26203 23545
rect 27154 23536 27160 23588
rect 27212 23576 27218 23588
rect 27212 23548 27752 23576
rect 27212 23536 27218 23548
rect 27724 23520 27752 23548
rect 30374 23536 30380 23588
rect 30432 23536 30438 23588
rect 18690 23508 18696 23520
rect 16776 23480 18696 23508
rect 18690 23468 18696 23480
rect 18748 23468 18754 23520
rect 19150 23468 19156 23520
rect 19208 23508 19214 23520
rect 22002 23508 22008 23520
rect 19208 23480 22008 23508
rect 19208 23468 19214 23480
rect 22002 23468 22008 23480
rect 22060 23468 22066 23520
rect 23106 23468 23112 23520
rect 23164 23508 23170 23520
rect 23293 23511 23351 23517
rect 23293 23508 23305 23511
rect 23164 23480 23305 23508
rect 23164 23468 23170 23480
rect 23293 23477 23305 23480
rect 23339 23477 23351 23511
rect 23293 23471 23351 23477
rect 27706 23468 27712 23520
rect 27764 23468 27770 23520
rect 28442 23468 28448 23520
rect 28500 23508 28506 23520
rect 30484 23508 30512 23675
rect 30558 23672 30564 23724
rect 30616 23712 30622 23724
rect 30926 23721 30932 23724
rect 30653 23715 30711 23721
rect 30653 23712 30665 23715
rect 30616 23684 30665 23712
rect 30616 23672 30622 23684
rect 30653 23681 30665 23684
rect 30699 23681 30711 23715
rect 30653 23675 30711 23681
rect 30883 23715 30932 23721
rect 30883 23681 30895 23715
rect 30929 23681 30932 23715
rect 30883 23675 30932 23681
rect 30668 23644 30696 23675
rect 30926 23672 30932 23675
rect 30984 23672 30990 23724
rect 30742 23644 30748 23656
rect 30668 23616 30748 23644
rect 30742 23604 30748 23616
rect 30800 23604 30806 23656
rect 28500 23480 30512 23508
rect 31021 23511 31079 23517
rect 28500 23468 28506 23480
rect 31021 23477 31033 23511
rect 31067 23508 31079 23511
rect 31662 23508 31668 23520
rect 31067 23480 31668 23508
rect 31067 23477 31079 23480
rect 31021 23471 31079 23477
rect 31662 23468 31668 23480
rect 31720 23468 31726 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 6730 23304 6736 23316
rect 6691 23276 6736 23304
rect 6730 23264 6736 23276
rect 6788 23264 6794 23316
rect 8205 23307 8263 23313
rect 8205 23273 8217 23307
rect 8251 23304 8263 23307
rect 8478 23304 8484 23316
rect 8251 23276 8484 23304
rect 8251 23273 8263 23276
rect 8205 23267 8263 23273
rect 8478 23264 8484 23276
rect 8536 23264 8542 23316
rect 10594 23264 10600 23316
rect 10652 23304 10658 23316
rect 10689 23307 10747 23313
rect 10689 23304 10701 23307
rect 10652 23276 10701 23304
rect 10652 23264 10658 23276
rect 10689 23273 10701 23276
rect 10735 23273 10747 23307
rect 10689 23267 10747 23273
rect 11241 23307 11299 23313
rect 11241 23273 11253 23307
rect 11287 23304 11299 23307
rect 11698 23304 11704 23316
rect 11287 23276 11704 23304
rect 11287 23273 11299 23276
rect 11241 23267 11299 23273
rect 11698 23264 11704 23276
rect 11756 23264 11762 23316
rect 13998 23264 14004 23316
rect 14056 23304 14062 23316
rect 14645 23307 14703 23313
rect 14645 23304 14657 23307
rect 14056 23276 14657 23304
rect 14056 23264 14062 23276
rect 14645 23273 14657 23276
rect 14691 23273 14703 23307
rect 14645 23267 14703 23273
rect 17037 23307 17095 23313
rect 17037 23273 17049 23307
rect 17083 23304 17095 23307
rect 17494 23304 17500 23316
rect 17083 23276 17500 23304
rect 17083 23273 17095 23276
rect 17037 23267 17095 23273
rect 17494 23264 17500 23276
rect 17552 23264 17558 23316
rect 18598 23304 18604 23316
rect 18559 23276 18604 23304
rect 18598 23264 18604 23276
rect 18656 23304 18662 23316
rect 20993 23307 21051 23313
rect 18656 23276 19334 23304
rect 18656 23264 18662 23276
rect 17218 23196 17224 23248
rect 17276 23236 17282 23248
rect 18874 23236 18880 23248
rect 17276 23208 18880 23236
rect 17276 23196 17282 23208
rect 18874 23196 18880 23208
rect 18932 23196 18938 23248
rect 19306 23236 19334 23276
rect 20993 23273 21005 23307
rect 21039 23304 21051 23307
rect 21174 23304 21180 23316
rect 21039 23276 21180 23304
rect 21039 23273 21051 23276
rect 20993 23267 21051 23273
rect 21174 23264 21180 23276
rect 21232 23264 21238 23316
rect 25498 23264 25504 23316
rect 25556 23304 25562 23316
rect 25593 23307 25651 23313
rect 25593 23304 25605 23307
rect 25556 23276 25605 23304
rect 25556 23264 25562 23276
rect 25593 23273 25605 23276
rect 25639 23273 25651 23307
rect 26234 23304 26240 23316
rect 26195 23276 26240 23304
rect 25593 23267 25651 23273
rect 26234 23264 26240 23276
rect 26292 23264 26298 23316
rect 28445 23307 28503 23313
rect 28445 23273 28457 23307
rect 28491 23304 28503 23307
rect 28718 23304 28724 23316
rect 28491 23276 28724 23304
rect 28491 23273 28503 23276
rect 28445 23267 28503 23273
rect 28718 23264 28724 23276
rect 28776 23264 28782 23316
rect 30006 23264 30012 23316
rect 30064 23304 30070 23316
rect 30558 23304 30564 23316
rect 30064 23276 30564 23304
rect 30064 23264 30070 23276
rect 30558 23264 30564 23276
rect 30616 23264 30622 23316
rect 22186 23236 22192 23248
rect 19306 23208 22192 23236
rect 22186 23196 22192 23208
rect 22244 23196 22250 23248
rect 8294 23128 8300 23180
rect 8352 23168 8358 23180
rect 8938 23168 8944 23180
rect 8352 23140 8944 23168
rect 8352 23128 8358 23140
rect 8938 23128 8944 23140
rect 8996 23168 9002 23180
rect 9309 23171 9367 23177
rect 9309 23168 9321 23171
rect 8996 23140 9321 23168
rect 8996 23128 9002 23140
rect 9309 23137 9321 23140
rect 9355 23137 9367 23171
rect 9309 23131 9367 23137
rect 16301 23171 16359 23177
rect 16301 23137 16313 23171
rect 16347 23168 16359 23171
rect 20714 23168 20720 23180
rect 16347 23140 17623 23168
rect 16347 23137 16359 23140
rect 16301 23131 16359 23137
rect 3786 23100 3792 23112
rect 3747 23072 3792 23100
rect 3786 23060 3792 23072
rect 3844 23060 3850 23112
rect 4056 23103 4114 23109
rect 4056 23069 4068 23103
rect 4102 23100 4114 23103
rect 4614 23100 4620 23112
rect 4102 23072 4620 23100
rect 4102 23069 4114 23072
rect 4056 23063 4114 23069
rect 4614 23060 4620 23072
rect 4672 23060 4678 23112
rect 6917 23103 6975 23109
rect 6917 23069 6929 23103
rect 6963 23100 6975 23103
rect 7282 23100 7288 23112
rect 6963 23072 7288 23100
rect 6963 23069 6975 23072
rect 6917 23063 6975 23069
rect 7282 23060 7288 23072
rect 7340 23060 7346 23112
rect 8389 23103 8447 23109
rect 8389 23069 8401 23103
rect 8435 23100 8447 23103
rect 9214 23100 9220 23112
rect 8435 23072 9220 23100
rect 8435 23069 8447 23072
rect 8389 23063 8447 23069
rect 9214 23060 9220 23072
rect 9272 23060 9278 23112
rect 11425 23103 11483 23109
rect 11425 23069 11437 23103
rect 11471 23100 11483 23103
rect 11790 23100 11796 23112
rect 11471 23072 11796 23100
rect 11471 23069 11483 23072
rect 11425 23063 11483 23069
rect 11790 23060 11796 23072
rect 11848 23060 11854 23112
rect 14277 23103 14335 23109
rect 14277 23069 14289 23103
rect 14323 23100 14335 23103
rect 14642 23100 14648 23112
rect 14323 23072 14648 23100
rect 14323 23069 14335 23072
rect 14277 23063 14335 23069
rect 14642 23060 14648 23072
rect 14700 23060 14706 23112
rect 16114 23100 16120 23112
rect 16027 23072 16120 23100
rect 16114 23060 16120 23072
rect 16172 23100 16178 23112
rect 16390 23100 16396 23112
rect 16172 23072 16396 23100
rect 16172 23060 16178 23072
rect 16390 23060 16396 23072
rect 16448 23060 16454 23112
rect 17218 23060 17224 23112
rect 17276 23109 17282 23112
rect 17276 23103 17325 23109
rect 17276 23069 17279 23103
rect 17313 23069 17325 23103
rect 17276 23063 17325 23069
rect 17405 23103 17463 23109
rect 17405 23069 17417 23103
rect 17451 23069 17463 23103
rect 17405 23063 17463 23069
rect 17497 23103 17555 23109
rect 17497 23069 17509 23103
rect 17543 23096 17555 23103
rect 17595 23096 17623 23140
rect 19628 23140 20720 23168
rect 17543 23069 17623 23096
rect 17497 23068 17623 23069
rect 17681 23103 17739 23109
rect 17681 23069 17693 23103
rect 17727 23100 17739 23103
rect 18322 23100 18328 23112
rect 17727 23072 18328 23100
rect 17727 23069 17739 23072
rect 17497 23063 17555 23068
rect 17681 23063 17739 23069
rect 17276 23060 17282 23063
rect 9576 23035 9634 23041
rect 9576 23001 9588 23035
rect 9622 23032 9634 23035
rect 10042 23032 10048 23044
rect 9622 23004 10048 23032
rect 9622 23001 9634 23004
rect 9576 22995 9634 23001
rect 10042 22992 10048 23004
rect 10100 22992 10106 23044
rect 13446 22992 13452 23044
rect 13504 23032 13510 23044
rect 14461 23035 14519 23041
rect 14461 23032 14473 23035
rect 13504 23004 14473 23032
rect 13504 22992 13510 23004
rect 14461 23001 14473 23004
rect 14507 23001 14519 23035
rect 14461 22995 14519 23001
rect 15933 23035 15991 23041
rect 15933 23001 15945 23035
rect 15979 23032 15991 23035
rect 16666 23032 16672 23044
rect 15979 23004 16672 23032
rect 15979 23001 15991 23004
rect 15933 22995 15991 23001
rect 16666 22992 16672 23004
rect 16724 22992 16730 23044
rect 17420 23032 17448 23063
rect 18322 23060 18328 23072
rect 18380 23060 18386 23112
rect 18417 23103 18475 23109
rect 18417 23069 18429 23103
rect 18463 23100 18475 23103
rect 18598 23100 18604 23112
rect 18463 23072 18604 23100
rect 18463 23069 18475 23072
rect 18417 23063 18475 23069
rect 18598 23060 18604 23072
rect 18656 23060 18662 23112
rect 19628 23032 19656 23140
rect 20714 23128 20720 23140
rect 20772 23168 20778 23180
rect 23750 23168 23756 23180
rect 20772 23140 23756 23168
rect 20772 23128 20778 23140
rect 19889 23103 19947 23109
rect 19889 23069 19901 23103
rect 19935 23100 19947 23103
rect 20254 23100 20260 23112
rect 19935 23072 20260 23100
rect 19935 23069 19947 23072
rect 19889 23063 19947 23069
rect 20254 23060 20260 23072
rect 20312 23100 20318 23112
rect 20806 23100 20812 23112
rect 20312 23072 20812 23100
rect 20312 23060 20318 23072
rect 20806 23060 20812 23072
rect 20864 23060 20870 23112
rect 22204 23109 22232 23140
rect 23750 23128 23756 23140
rect 23808 23128 23814 23180
rect 25240 23140 28120 23168
rect 22097 23103 22155 23109
rect 22097 23069 22109 23103
rect 22143 23069 22155 23103
rect 22097 23063 22155 23069
rect 22189 23103 22247 23109
rect 22189 23069 22201 23103
rect 22235 23069 22247 23103
rect 22189 23063 22247 23069
rect 17420 23004 19656 23032
rect 19705 23035 19763 23041
rect 19705 23001 19717 23035
rect 19751 23032 19763 23035
rect 20349 23035 20407 23041
rect 20349 23032 20361 23035
rect 19751 23004 20361 23032
rect 19751 23001 19763 23004
rect 19705 22995 19763 23001
rect 20349 23001 20361 23004
rect 20395 23001 20407 23035
rect 20898 23032 20904 23044
rect 20859 23004 20904 23032
rect 20349 22995 20407 23001
rect 4706 22924 4712 22976
rect 4764 22964 4770 22976
rect 5169 22967 5227 22973
rect 5169 22964 5181 22967
rect 4764 22936 5181 22964
rect 4764 22924 4770 22936
rect 5169 22933 5181 22936
rect 5215 22933 5227 22967
rect 5169 22927 5227 22933
rect 12342 22924 12348 22976
rect 12400 22964 12406 22976
rect 19720 22964 19748 22995
rect 12400 22936 19748 22964
rect 20073 22967 20131 22973
rect 12400 22924 12406 22936
rect 20073 22933 20085 22967
rect 20119 22964 20131 22967
rect 20254 22964 20260 22976
rect 20119 22936 20260 22964
rect 20119 22933 20131 22936
rect 20073 22927 20131 22933
rect 20254 22924 20260 22936
rect 20312 22924 20318 22976
rect 20364 22964 20392 22995
rect 20898 22992 20904 23004
rect 20956 22992 20962 23044
rect 22112 23032 22140 23063
rect 22278 23060 22284 23112
rect 22336 23100 22342 23112
rect 22465 23103 22523 23109
rect 22336 23072 22381 23100
rect 22336 23060 22342 23072
rect 22465 23069 22477 23103
rect 22511 23100 22523 23103
rect 22554 23100 22560 23112
rect 22511 23072 22560 23100
rect 22511 23069 22523 23072
rect 22465 23063 22523 23069
rect 22554 23060 22560 23072
rect 22612 23100 22618 23112
rect 23382 23100 23388 23112
rect 22612 23072 23388 23100
rect 22612 23060 22618 23072
rect 23382 23060 23388 23072
rect 23440 23060 23446 23112
rect 25038 23060 25044 23112
rect 25096 23100 25102 23112
rect 25240 23109 25268 23140
rect 25225 23103 25283 23109
rect 25225 23100 25237 23103
rect 25096 23072 25237 23100
rect 25096 23060 25102 23072
rect 25225 23069 25237 23072
rect 25271 23069 25283 23103
rect 25225 23063 25283 23069
rect 25409 23103 25467 23109
rect 25409 23069 25421 23103
rect 25455 23100 25467 23103
rect 26418 23100 26424 23112
rect 25455 23072 26424 23100
rect 25455 23069 25467 23072
rect 25409 23063 25467 23069
rect 26418 23060 26424 23072
rect 26476 23060 26482 23112
rect 28092 23109 28120 23140
rect 28077 23103 28135 23109
rect 28077 23069 28089 23103
rect 28123 23069 28135 23103
rect 28077 23063 28135 23069
rect 28261 23103 28319 23109
rect 28261 23069 28273 23103
rect 28307 23100 28319 23103
rect 28442 23100 28448 23112
rect 28307 23072 28448 23100
rect 28307 23069 28319 23072
rect 28261 23063 28319 23069
rect 28442 23060 28448 23072
rect 28500 23060 28506 23112
rect 32674 23100 32680 23112
rect 32635 23072 32680 23100
rect 32674 23060 32680 23072
rect 32732 23060 32738 23112
rect 23474 23032 23480 23044
rect 22112 23004 23480 23032
rect 23474 22992 23480 23004
rect 23532 22992 23538 23044
rect 25774 22992 25780 23044
rect 25832 23032 25838 23044
rect 26145 23035 26203 23041
rect 26145 23032 26157 23035
rect 25832 23004 26157 23032
rect 25832 22992 25838 23004
rect 26145 23001 26157 23004
rect 26191 23001 26203 23035
rect 26145 22995 26203 23001
rect 21174 22964 21180 22976
rect 20364 22936 21180 22964
rect 21174 22924 21180 22936
rect 21232 22924 21238 22976
rect 21821 22967 21879 22973
rect 21821 22933 21833 22967
rect 21867 22964 21879 22967
rect 21910 22964 21916 22976
rect 21867 22936 21916 22964
rect 21867 22933 21879 22936
rect 21821 22927 21879 22933
rect 21910 22924 21916 22936
rect 21968 22924 21974 22976
rect 22186 22924 22192 22976
rect 22244 22964 22250 22976
rect 22554 22964 22560 22976
rect 22244 22936 22560 22964
rect 22244 22924 22250 22936
rect 22554 22924 22560 22936
rect 22612 22924 22618 22976
rect 32490 22964 32496 22976
rect 32451 22936 32496 22964
rect 32490 22924 32496 22936
rect 32548 22924 32554 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 2746 22732 12434 22760
rect 14 22516 20 22568
rect 72 22556 78 22568
rect 2746 22556 2774 22732
rect 4525 22695 4583 22701
rect 4525 22661 4537 22695
rect 4571 22661 4583 22695
rect 4525 22655 4583 22661
rect 4741 22695 4799 22701
rect 4741 22661 4753 22695
rect 4787 22692 4799 22695
rect 5442 22692 5448 22704
rect 4787 22664 5448 22692
rect 4787 22661 4799 22664
rect 4741 22655 4799 22661
rect 4540 22624 4568 22655
rect 5442 22652 5448 22664
rect 5500 22652 5506 22704
rect 6549 22695 6607 22701
rect 6549 22661 6561 22695
rect 6595 22661 6607 22695
rect 6549 22655 6607 22661
rect 6765 22695 6823 22701
rect 6765 22661 6777 22695
rect 6811 22692 6823 22695
rect 7834 22692 7840 22704
rect 6811 22664 7840 22692
rect 6811 22661 6823 22664
rect 6765 22655 6823 22661
rect 5718 22624 5724 22636
rect 4540 22596 5724 22624
rect 5718 22584 5724 22596
rect 5776 22584 5782 22636
rect 72 22528 2774 22556
rect 6564 22556 6592 22655
rect 7834 22652 7840 22664
rect 7892 22652 7898 22704
rect 11514 22692 11520 22704
rect 11475 22664 11520 22692
rect 11514 22652 11520 22664
rect 11572 22652 11578 22704
rect 11698 22652 11704 22704
rect 11756 22701 11762 22704
rect 11756 22695 11775 22701
rect 11763 22661 11775 22695
rect 12406 22692 12434 22732
rect 13446 22720 13452 22772
rect 13504 22760 13510 22772
rect 14369 22763 14427 22769
rect 14369 22760 14381 22763
rect 13504 22732 14381 22760
rect 13504 22720 13510 22732
rect 14369 22729 14381 22732
rect 14415 22729 14427 22763
rect 14369 22723 14427 22729
rect 18138 22720 18144 22772
rect 18196 22760 18202 22772
rect 19978 22760 19984 22772
rect 18196 22732 19984 22760
rect 18196 22720 18202 22732
rect 19978 22720 19984 22732
rect 20036 22760 20042 22772
rect 20717 22763 20775 22769
rect 20717 22760 20729 22763
rect 20036 22732 20729 22760
rect 20036 22720 20042 22732
rect 20717 22729 20729 22732
rect 20763 22729 20775 22763
rect 20717 22723 20775 22729
rect 23201 22763 23259 22769
rect 23201 22729 23213 22763
rect 23247 22760 23259 22763
rect 23474 22760 23480 22772
rect 23247 22732 23480 22760
rect 23247 22729 23259 22732
rect 23201 22723 23259 22729
rect 23474 22720 23480 22732
rect 23532 22720 23538 22772
rect 23753 22763 23811 22769
rect 23753 22729 23765 22763
rect 23799 22760 23811 22763
rect 23934 22760 23940 22772
rect 23799 22732 23940 22760
rect 23799 22729 23811 22732
rect 23753 22723 23811 22729
rect 23934 22720 23940 22732
rect 23992 22720 23998 22772
rect 26418 22760 26424 22772
rect 26379 22732 26424 22760
rect 26418 22720 26424 22732
rect 26476 22720 26482 22772
rect 19429 22695 19487 22701
rect 19429 22692 19441 22695
rect 12406 22664 19441 22692
rect 11756 22655 11775 22661
rect 19429 22661 19441 22664
rect 19475 22661 19487 22695
rect 22462 22692 22468 22704
rect 19429 22655 19487 22661
rect 21836 22664 22468 22692
rect 11756 22652 11762 22655
rect 7190 22584 7196 22636
rect 7248 22624 7254 22636
rect 7561 22627 7619 22633
rect 7561 22624 7573 22627
rect 7248 22596 7573 22624
rect 7248 22584 7254 22596
rect 7561 22593 7573 22596
rect 7607 22593 7619 22627
rect 7561 22587 7619 22593
rect 8297 22627 8355 22633
rect 8297 22593 8309 22627
rect 8343 22624 8355 22627
rect 8662 22624 8668 22636
rect 8343 22596 8668 22624
rect 8343 22593 8355 22596
rect 8297 22587 8355 22593
rect 8662 22584 8668 22596
rect 8720 22584 8726 22636
rect 10229 22627 10287 22633
rect 10229 22593 10241 22627
rect 10275 22624 10287 22627
rect 10778 22624 10784 22636
rect 10275 22596 10784 22624
rect 10275 22593 10287 22596
rect 10229 22587 10287 22593
rect 10778 22584 10784 22596
rect 10836 22584 10842 22636
rect 11238 22584 11244 22636
rect 11296 22624 11302 22636
rect 11716 22624 11744 22652
rect 11296 22596 11744 22624
rect 12529 22627 12587 22633
rect 11296 22584 11302 22596
rect 12529 22593 12541 22627
rect 12575 22624 12587 22627
rect 12894 22624 12900 22636
rect 12575 22596 12900 22624
rect 12575 22593 12587 22596
rect 12529 22587 12587 22593
rect 12894 22584 12900 22596
rect 12952 22584 12958 22636
rect 13078 22584 13084 22636
rect 13136 22624 13142 22636
rect 13245 22627 13303 22633
rect 13245 22624 13257 22627
rect 13136 22596 13257 22624
rect 13136 22584 13142 22596
rect 13245 22593 13257 22596
rect 13291 22593 13303 22627
rect 13245 22587 13303 22593
rect 17497 22627 17555 22633
rect 17497 22593 17509 22627
rect 17543 22624 17555 22627
rect 18230 22624 18236 22636
rect 17543 22596 18236 22624
rect 17543 22593 17555 22596
rect 17497 22587 17555 22593
rect 18230 22584 18236 22596
rect 18288 22584 18294 22636
rect 18325 22627 18383 22633
rect 18325 22593 18337 22627
rect 18371 22624 18383 22627
rect 19242 22624 19248 22636
rect 18371 22596 19248 22624
rect 18371 22593 18383 22596
rect 18325 22587 18383 22593
rect 19242 22584 19248 22596
rect 19300 22584 19306 22636
rect 21836 22633 21864 22664
rect 22462 22652 22468 22664
rect 22520 22692 22526 22704
rect 29270 22692 29276 22704
rect 22520 22664 25084 22692
rect 22520 22652 22526 22664
rect 25056 22636 25084 22664
rect 27724 22664 29276 22692
rect 21821 22627 21879 22633
rect 21821 22593 21833 22627
rect 21867 22593 21879 22627
rect 21821 22587 21879 22593
rect 21910 22584 21916 22636
rect 21968 22624 21974 22636
rect 22077 22627 22135 22633
rect 22077 22624 22089 22627
rect 21968 22596 22089 22624
rect 21968 22584 21974 22596
rect 22077 22593 22089 22596
rect 22123 22593 22135 22627
rect 22077 22587 22135 22593
rect 23474 22584 23480 22636
rect 23532 22624 23538 22636
rect 23661 22627 23719 22633
rect 23661 22624 23673 22627
rect 23532 22596 23673 22624
rect 23532 22584 23538 22596
rect 23661 22593 23673 22596
rect 23707 22593 23719 22627
rect 23842 22624 23848 22636
rect 23803 22596 23848 22624
rect 23661 22587 23719 22593
rect 8570 22556 8576 22568
rect 6564 22528 7420 22556
rect 8531 22528 8576 22556
rect 72 22516 78 22528
rect 7392 22500 7420 22528
rect 8570 22516 8576 22528
rect 8628 22516 8634 22568
rect 12434 22516 12440 22568
rect 12492 22556 12498 22568
rect 12989 22559 13047 22565
rect 12989 22556 13001 22559
rect 12492 22528 13001 22556
rect 12492 22516 12498 22528
rect 12989 22525 13001 22528
rect 13035 22525 13047 22559
rect 12989 22519 13047 22525
rect 18141 22559 18199 22565
rect 18141 22525 18153 22559
rect 18187 22556 18199 22559
rect 18782 22556 18788 22568
rect 18187 22528 18788 22556
rect 18187 22525 18199 22528
rect 18141 22519 18199 22525
rect 18782 22516 18788 22528
rect 18840 22516 18846 22568
rect 23676 22556 23704 22587
rect 23842 22584 23848 22596
rect 23900 22584 23906 22636
rect 25038 22624 25044 22636
rect 24951 22596 25044 22624
rect 25038 22584 25044 22596
rect 25096 22584 25102 22636
rect 25130 22584 25136 22636
rect 25188 22624 25194 22636
rect 27724 22633 27752 22664
rect 29270 22652 29276 22664
rect 29328 22652 29334 22704
rect 30558 22692 30564 22704
rect 30208 22664 30564 22692
rect 25297 22627 25355 22633
rect 25297 22624 25309 22627
rect 25188 22596 25309 22624
rect 25188 22584 25194 22596
rect 25297 22593 25309 22596
rect 25343 22593 25355 22627
rect 25297 22587 25355 22593
rect 27709 22627 27767 22633
rect 27709 22593 27721 22627
rect 27755 22593 27767 22627
rect 27801 22627 27859 22633
rect 27801 22624 27813 22627
rect 27709 22587 27767 22593
rect 27797 22593 27813 22624
rect 27847 22593 27859 22627
rect 27797 22587 27859 22593
rect 23750 22556 23756 22568
rect 23676 22528 23756 22556
rect 23750 22516 23756 22528
rect 23808 22516 23814 22568
rect 27338 22516 27344 22568
rect 27396 22556 27402 22568
rect 27797 22556 27825 22587
rect 27890 22584 27896 22636
rect 27948 22624 27954 22636
rect 28077 22627 28135 22633
rect 27948 22596 27993 22624
rect 27948 22584 27954 22596
rect 28077 22593 28089 22627
rect 28123 22624 28135 22627
rect 28350 22624 28356 22636
rect 28123 22596 28356 22624
rect 28123 22593 28135 22596
rect 28077 22587 28135 22593
rect 28350 22584 28356 22596
rect 28408 22584 28414 22636
rect 29914 22584 29920 22636
rect 29972 22624 29978 22636
rect 30208 22633 30236 22664
rect 30558 22652 30564 22664
rect 30616 22692 30622 22704
rect 32392 22695 32450 22701
rect 30616 22664 32168 22692
rect 30616 22652 30622 22664
rect 30193 22627 30251 22633
rect 30193 22624 30205 22627
rect 29972 22596 30205 22624
rect 29972 22584 29978 22596
rect 30193 22593 30205 22596
rect 30239 22593 30251 22627
rect 30193 22587 30251 22593
rect 30460 22627 30518 22633
rect 30460 22593 30472 22627
rect 30506 22624 30518 22627
rect 30926 22624 30932 22636
rect 30506 22596 30932 22624
rect 30506 22593 30518 22596
rect 30460 22587 30518 22593
rect 30926 22584 30932 22596
rect 30984 22584 30990 22636
rect 32140 22633 32168 22664
rect 32392 22661 32404 22695
rect 32438 22692 32450 22695
rect 32490 22692 32496 22704
rect 32438 22664 32496 22692
rect 32438 22661 32450 22664
rect 32392 22655 32450 22661
rect 32490 22652 32496 22664
rect 32548 22652 32554 22704
rect 32125 22627 32183 22633
rect 32125 22593 32137 22627
rect 32171 22593 32183 22627
rect 34146 22624 34152 22636
rect 34107 22596 34152 22624
rect 32125 22587 32183 22593
rect 34146 22584 34152 22596
rect 34204 22584 34210 22636
rect 27396 22528 27825 22556
rect 27396 22516 27402 22528
rect 4890 22488 4896 22500
rect 4851 22460 4896 22488
rect 4890 22448 4896 22460
rect 4948 22448 4954 22500
rect 7006 22488 7012 22500
rect 6748 22460 7012 22488
rect 4706 22420 4712 22432
rect 4667 22392 4712 22420
rect 4706 22380 4712 22392
rect 4764 22380 4770 22432
rect 6748 22429 6776 22460
rect 7006 22448 7012 22460
rect 7064 22448 7070 22500
rect 7374 22488 7380 22500
rect 7335 22460 7380 22488
rect 7374 22448 7380 22460
rect 7432 22448 7438 22500
rect 10042 22488 10048 22500
rect 10003 22460 10048 22488
rect 10042 22448 10048 22460
rect 10100 22448 10106 22500
rect 12158 22488 12164 22500
rect 11716 22460 12164 22488
rect 6733 22423 6791 22429
rect 6733 22389 6745 22423
rect 6779 22389 6791 22423
rect 6914 22420 6920 22432
rect 6875 22392 6920 22420
rect 6733 22383 6791 22389
rect 6914 22380 6920 22392
rect 6972 22380 6978 22432
rect 11716 22429 11744 22460
rect 12158 22448 12164 22460
rect 12216 22448 12222 22500
rect 17770 22448 17776 22500
rect 17828 22488 17834 22500
rect 20714 22488 20720 22500
rect 17828 22460 20720 22488
rect 17828 22448 17834 22460
rect 20714 22448 20720 22460
rect 20772 22448 20778 22500
rect 11701 22423 11759 22429
rect 11701 22389 11713 22423
rect 11747 22389 11759 22423
rect 11882 22420 11888 22432
rect 11843 22392 11888 22420
rect 11701 22383 11759 22389
rect 11882 22380 11888 22392
rect 11940 22380 11946 22432
rect 12342 22420 12348 22432
rect 12303 22392 12348 22420
rect 12342 22380 12348 22392
rect 12400 22380 12406 22432
rect 17494 22380 17500 22432
rect 17552 22420 17558 22432
rect 17589 22423 17647 22429
rect 17589 22420 17601 22423
rect 17552 22392 17601 22420
rect 17552 22380 17558 22392
rect 17589 22389 17601 22392
rect 17635 22389 17647 22423
rect 17589 22383 17647 22389
rect 18138 22380 18144 22432
rect 18196 22420 18202 22432
rect 18509 22423 18567 22429
rect 18509 22420 18521 22423
rect 18196 22392 18521 22420
rect 18196 22380 18202 22392
rect 18509 22389 18521 22392
rect 18555 22389 18567 22423
rect 18509 22383 18567 22389
rect 27433 22423 27491 22429
rect 27433 22389 27445 22423
rect 27479 22420 27491 22423
rect 27706 22420 27712 22432
rect 27479 22392 27712 22420
rect 27479 22389 27491 22392
rect 27433 22383 27491 22389
rect 27706 22380 27712 22392
rect 27764 22380 27770 22432
rect 28074 22380 28080 22432
rect 28132 22420 28138 22432
rect 28902 22420 28908 22432
rect 28132 22392 28908 22420
rect 28132 22380 28138 22392
rect 28902 22380 28908 22392
rect 28960 22380 28966 22432
rect 31294 22380 31300 22432
rect 31352 22420 31358 22432
rect 31573 22423 31631 22429
rect 31573 22420 31585 22423
rect 31352 22392 31585 22420
rect 31352 22380 31358 22392
rect 31573 22389 31585 22392
rect 31619 22389 31631 22423
rect 33502 22420 33508 22432
rect 33463 22392 33508 22420
rect 31573 22383 31631 22389
rect 33502 22380 33508 22392
rect 33560 22380 33566 22432
rect 33962 22420 33968 22432
rect 33923 22392 33968 22420
rect 33962 22380 33968 22392
rect 34020 22380 34026 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 7006 22216 7012 22228
rect 6967 22188 7012 22216
rect 7006 22176 7012 22188
rect 7064 22176 7070 22228
rect 8662 22176 8668 22228
rect 8720 22216 8726 22228
rect 12158 22216 12164 22228
rect 8720 22188 11744 22216
rect 12119 22188 12164 22216
rect 8720 22176 8726 22188
rect 11716 22148 11744 22188
rect 12158 22176 12164 22188
rect 12216 22176 12222 22228
rect 12802 22216 12808 22228
rect 12763 22188 12808 22216
rect 12802 22176 12808 22188
rect 12860 22176 12866 22228
rect 12894 22176 12900 22228
rect 12952 22216 12958 22228
rect 13078 22216 13084 22228
rect 12952 22188 13084 22216
rect 12952 22176 12958 22188
rect 13078 22176 13084 22188
rect 13136 22176 13142 22228
rect 14660 22188 18184 22216
rect 14660 22148 14688 22188
rect 11716 22120 14688 22148
rect 18156 22148 18184 22188
rect 18230 22176 18236 22228
rect 18288 22216 18294 22228
rect 18509 22219 18567 22225
rect 18509 22216 18521 22219
rect 18288 22188 18521 22216
rect 18288 22176 18294 22188
rect 18509 22185 18521 22188
rect 18555 22216 18567 22219
rect 19150 22216 19156 22228
rect 18555 22188 19156 22216
rect 18555 22185 18567 22188
rect 18509 22179 18567 22185
rect 19150 22176 19156 22188
rect 19208 22176 19214 22228
rect 20898 22216 20904 22228
rect 19812 22188 20904 22216
rect 19812 22148 19840 22188
rect 20898 22176 20904 22188
rect 20956 22216 20962 22228
rect 21542 22216 21548 22228
rect 20956 22188 21548 22216
rect 20956 22176 20962 22188
rect 21542 22176 21548 22188
rect 21600 22176 21606 22228
rect 28442 22216 28448 22228
rect 27448 22188 28448 22216
rect 18156 22120 19840 22148
rect 20806 22108 20812 22160
rect 20864 22148 20870 22160
rect 21177 22151 21235 22157
rect 21177 22148 21189 22151
rect 20864 22120 21189 22148
rect 20864 22108 20870 22120
rect 21177 22117 21189 22120
rect 21223 22117 21235 22151
rect 25774 22148 25780 22160
rect 21177 22111 21235 22117
rect 25516 22120 25780 22148
rect 5442 22040 5448 22092
rect 5500 22080 5506 22092
rect 7469 22083 7527 22089
rect 5500 22052 5764 22080
rect 5500 22040 5506 22052
rect 3786 21972 3792 22024
rect 3844 22012 3850 22024
rect 5629 22015 5687 22021
rect 5629 22012 5641 22015
rect 3844 21984 5641 22012
rect 3844 21972 3850 21984
rect 5629 21981 5641 21984
rect 5675 21981 5687 22015
rect 5736 22012 5764 22052
rect 7469 22049 7481 22083
rect 7515 22080 7527 22083
rect 8662 22080 8668 22092
rect 7515 22052 8668 22080
rect 7515 22049 7527 22052
rect 7469 22043 7527 22049
rect 8662 22040 8668 22052
rect 8720 22040 8726 22092
rect 12894 22040 12900 22092
rect 12952 22080 12958 22092
rect 12952 22052 14780 22080
rect 12952 22040 12958 22052
rect 7745 22015 7803 22021
rect 7745 22012 7757 22015
rect 5736 21984 7757 22012
rect 5629 21975 5687 21981
rect 7745 21981 7757 21984
rect 7791 21981 7803 22015
rect 7745 21975 7803 21981
rect 10781 22015 10839 22021
rect 10781 21981 10793 22015
rect 10827 22012 10839 22015
rect 10870 22012 10876 22024
rect 10827 21984 10876 22012
rect 10827 21981 10839 21984
rect 10781 21975 10839 21981
rect 10870 21972 10876 21984
rect 10928 22012 10934 22024
rect 12434 22012 12440 22024
rect 10928 21984 12440 22012
rect 10928 21972 10934 21984
rect 12434 21972 12440 21984
rect 12492 21972 12498 22024
rect 14090 21972 14096 22024
rect 14148 22012 14154 22024
rect 14645 22015 14703 22021
rect 14645 22012 14657 22015
rect 14148 21984 14657 22012
rect 14148 21972 14154 21984
rect 14645 21981 14657 21984
rect 14691 21981 14703 22015
rect 14752 22012 14780 22052
rect 17954 22040 17960 22092
rect 18012 22080 18018 22092
rect 22462 22080 22468 22092
rect 18012 22052 19932 22080
rect 22423 22052 22468 22080
rect 18012 22040 18018 22052
rect 15654 22012 15660 22024
rect 14752 21984 15660 22012
rect 14645 21975 14703 21981
rect 15654 21972 15660 21984
rect 15712 21972 15718 22024
rect 16485 22015 16543 22021
rect 16485 21981 16497 22015
rect 16531 22012 16543 22015
rect 17310 22012 17316 22024
rect 16531 21984 17316 22012
rect 16531 21981 16543 21984
rect 16485 21975 16543 21981
rect 17310 21972 17316 21984
rect 17368 22012 17374 22024
rect 19797 22015 19855 22021
rect 19797 22012 19809 22015
rect 17368 21984 19809 22012
rect 17368 21972 17374 21984
rect 19797 21981 19809 21984
rect 19843 21981 19855 22015
rect 19904 22012 19932 22052
rect 22462 22040 22468 22052
rect 22520 22040 22526 22092
rect 23934 22040 23940 22092
rect 23992 22080 23998 22092
rect 25516 22080 25544 22120
rect 23992 22052 25544 22080
rect 23992 22040 23998 22052
rect 24596 22021 24624 22052
rect 24762 22021 24768 22024
rect 24581 22015 24639 22021
rect 19904 21984 24440 22012
rect 19797 21975 19855 21981
rect 5896 21947 5954 21953
rect 5896 21913 5908 21947
rect 5942 21944 5954 21947
rect 6270 21944 6276 21956
rect 5942 21916 6276 21944
rect 5942 21913 5954 21916
rect 5896 21907 5954 21913
rect 6270 21904 6276 21916
rect 6328 21904 6334 21956
rect 11048 21947 11106 21953
rect 11048 21913 11060 21947
rect 11094 21944 11106 21947
rect 11330 21944 11336 21956
rect 11094 21916 11336 21944
rect 11094 21913 11106 21916
rect 11048 21907 11106 21913
rect 11330 21904 11336 21916
rect 11388 21904 11394 21956
rect 11514 21904 11520 21956
rect 11572 21944 11578 21956
rect 12621 21947 12679 21953
rect 12621 21944 12633 21947
rect 11572 21916 12633 21944
rect 11572 21904 11578 21916
rect 12621 21913 12633 21916
rect 12667 21913 12679 21947
rect 12621 21907 12679 21913
rect 14912 21947 14970 21953
rect 14912 21913 14924 21947
rect 14958 21944 14970 21947
rect 15562 21944 15568 21956
rect 14958 21916 15568 21944
rect 14958 21913 14970 21916
rect 14912 21907 14970 21913
rect 15562 21904 15568 21916
rect 15620 21904 15626 21956
rect 16206 21904 16212 21956
rect 16264 21944 16270 21956
rect 16730 21947 16788 21953
rect 16730 21944 16742 21947
rect 16264 21916 16742 21944
rect 16264 21904 16270 21916
rect 16730 21913 16742 21916
rect 16776 21913 16788 21947
rect 16730 21907 16788 21913
rect 18325 21947 18383 21953
rect 18325 21913 18337 21947
rect 18371 21944 18383 21947
rect 19058 21944 19064 21956
rect 18371 21916 19064 21944
rect 18371 21913 18383 21916
rect 18325 21907 18383 21913
rect 19058 21904 19064 21916
rect 19116 21904 19122 21956
rect 20070 21953 20076 21956
rect 20064 21907 20076 21953
rect 20128 21944 20134 21956
rect 21821 21947 21879 21953
rect 20128 21916 20164 21944
rect 20070 21904 20076 21907
rect 20128 21904 20134 21916
rect 21821 21913 21833 21947
rect 21867 21944 21879 21947
rect 22094 21944 22100 21956
rect 21867 21916 22100 21944
rect 21867 21913 21879 21916
rect 21821 21907 21879 21913
rect 22094 21904 22100 21916
rect 22152 21904 22158 21956
rect 22732 21947 22790 21953
rect 22732 21913 22744 21947
rect 22778 21944 22790 21947
rect 22830 21944 22836 21956
rect 22778 21916 22836 21944
rect 22778 21913 22790 21916
rect 22732 21907 22790 21913
rect 22830 21904 22836 21916
rect 22888 21904 22894 21956
rect 24412 21944 24440 21984
rect 24581 21981 24593 22015
rect 24627 21981 24639 22015
rect 24581 21975 24639 21981
rect 24729 22015 24768 22021
rect 24729 21981 24741 22015
rect 24729 21975 24768 21981
rect 24762 21972 24768 21975
rect 24820 21972 24826 22024
rect 24946 22012 24952 22024
rect 24907 21984 24952 22012
rect 24946 21972 24952 21984
rect 25004 21972 25010 22024
rect 25130 22021 25136 22024
rect 25087 22015 25136 22021
rect 25087 21981 25099 22015
rect 25133 21981 25136 22015
rect 25087 21975 25136 21981
rect 25130 21972 25136 21975
rect 25188 21972 25194 22024
rect 25700 22021 25728 22120
rect 25774 22108 25780 22120
rect 25832 22108 25838 22160
rect 26418 22148 26424 22160
rect 25884 22120 26424 22148
rect 25884 22021 25912 22120
rect 26418 22108 26424 22120
rect 26476 22108 26482 22160
rect 26510 22040 26516 22092
rect 26568 22080 26574 22092
rect 27448 22080 27476 22188
rect 28442 22176 28448 22188
rect 28500 22176 28506 22228
rect 28813 22219 28871 22225
rect 28813 22185 28825 22219
rect 28859 22216 28871 22219
rect 28902 22216 28908 22228
rect 28859 22188 28908 22216
rect 28859 22185 28871 22188
rect 28813 22179 28871 22185
rect 28902 22176 28908 22188
rect 28960 22176 28966 22228
rect 30926 22216 30932 22228
rect 30887 22188 30932 22216
rect 30926 22176 30932 22188
rect 30984 22176 30990 22228
rect 30098 22108 30104 22160
rect 30156 22108 30162 22160
rect 30190 22108 30196 22160
rect 30248 22108 30254 22160
rect 29822 22080 29828 22092
rect 26568 22052 27476 22080
rect 29783 22052 29828 22080
rect 26568 22040 26574 22052
rect 29822 22040 29828 22052
rect 29880 22040 29886 22092
rect 25685 22015 25743 22021
rect 25685 21981 25697 22015
rect 25731 21981 25743 22015
rect 25685 21975 25743 21981
rect 25833 22015 25912 22021
rect 25833 21981 25845 22015
rect 25879 21984 25912 22015
rect 26050 22012 26056 22024
rect 26011 21984 26056 22012
rect 25879 21981 25891 21984
rect 25833 21975 25891 21981
rect 26050 21972 26056 21984
rect 26108 21972 26114 22024
rect 26142 21972 26148 22024
rect 26200 22021 26206 22024
rect 26200 22012 26208 22021
rect 26602 22012 26608 22024
rect 26200 21984 26608 22012
rect 26200 21975 26208 21984
rect 26200 21972 26206 21975
rect 26602 21972 26608 21984
rect 26660 21972 26666 22024
rect 27433 22015 27491 22021
rect 27433 21981 27445 22015
rect 27479 22012 27491 22015
rect 27479 21984 28212 22012
rect 27479 21981 27491 21984
rect 27433 21975 27491 21981
rect 24857 21947 24915 21953
rect 24857 21944 24869 21947
rect 24412 21916 24869 21944
rect 24857 21913 24869 21916
rect 24903 21944 24915 21947
rect 25961 21947 26019 21953
rect 25961 21944 25973 21947
rect 24903 21916 25973 21944
rect 24903 21913 24915 21916
rect 24857 21907 24915 21913
rect 25792 21888 25820 21916
rect 25961 21913 25973 21916
rect 26007 21913 26019 21947
rect 25961 21907 26019 21913
rect 27686 21904 27692 21956
rect 27744 21944 27750 21956
rect 28184 21944 28212 21984
rect 28810 21972 28816 22024
rect 28868 22012 28874 22024
rect 30116 22021 30144 22108
rect 30209 22080 30237 22108
rect 30742 22080 30748 22092
rect 30209 22052 30333 22080
rect 30305 22021 30333 22052
rect 30484 22052 30748 22080
rect 30484 22024 30512 22052
rect 30742 22040 30748 22052
rect 30800 22080 30806 22092
rect 32953 22083 33011 22089
rect 30800 22052 31616 22080
rect 30800 22040 30806 22052
rect 30101 22015 30159 22021
rect 28868 21984 30052 22012
rect 28868 21972 28874 21984
rect 29914 21944 29920 21956
rect 27744 21916 27789 21944
rect 28184 21916 29920 21944
rect 27744 21904 27750 21916
rect 29914 21904 29920 21916
rect 29972 21904 29978 21956
rect 30024 21944 30052 21984
rect 30101 21981 30113 22015
rect 30147 21981 30159 22015
rect 30101 21975 30159 21981
rect 30193 22015 30251 22021
rect 30193 21981 30205 22015
rect 30239 21981 30251 22015
rect 30193 21975 30251 21981
rect 30290 22015 30348 22021
rect 30290 21981 30302 22015
rect 30336 21981 30348 22015
rect 30290 21975 30348 21981
rect 30208 21944 30236 21975
rect 30466 21972 30472 22024
rect 30524 22012 30530 22024
rect 30524 21984 30569 22012
rect 30524 21972 30530 21984
rect 30834 21972 30840 22024
rect 30892 22012 30898 22024
rect 31202 22012 31208 22024
rect 30892 21984 31208 22012
rect 30892 21972 30898 21984
rect 31202 21972 31208 21984
rect 31260 21972 31266 22024
rect 31297 22015 31355 22021
rect 31297 21981 31309 22015
rect 31343 21981 31355 22015
rect 31297 21975 31355 21981
rect 30650 21944 30656 21956
rect 30024 21916 30656 21944
rect 30650 21904 30656 21916
rect 30708 21944 30714 21956
rect 31312 21944 31340 21975
rect 31386 21972 31392 22024
rect 31444 22012 31450 22024
rect 31588 22021 31616 22052
rect 32953 22049 32965 22083
rect 32999 22080 33011 22083
rect 33502 22080 33508 22092
rect 32999 22052 33508 22080
rect 32999 22049 33011 22052
rect 32953 22043 33011 22049
rect 33502 22040 33508 22052
rect 33560 22040 33566 22092
rect 34057 22083 34115 22089
rect 34057 22080 34069 22083
rect 33612 22052 34069 22080
rect 31573 22015 31631 22021
rect 31444 21984 31489 22012
rect 31444 21972 31450 21984
rect 31573 21981 31585 22015
rect 31619 21981 31631 22015
rect 31573 21975 31631 21981
rect 31662 21972 31668 22024
rect 31720 22012 31726 22024
rect 32677 22015 32735 22021
rect 32677 22012 32689 22015
rect 31720 21984 32689 22012
rect 31720 21972 31726 21984
rect 32677 21981 32689 21984
rect 32723 21981 32735 22015
rect 32677 21975 32735 21981
rect 32858 21972 32864 22024
rect 32916 22012 32922 22024
rect 33612 22012 33640 22052
rect 34057 22049 34069 22052
rect 34103 22049 34115 22083
rect 34057 22043 34115 22049
rect 32916 21984 33640 22012
rect 33873 22015 33931 22021
rect 32916 21972 32922 21984
rect 33873 21981 33885 22015
rect 33919 21981 33931 22015
rect 33873 21975 33931 21981
rect 34149 22015 34207 22021
rect 34149 21981 34161 22015
rect 34195 22012 34207 22015
rect 34974 22012 34980 22024
rect 34195 21984 34980 22012
rect 34195 21981 34207 21984
rect 34149 21975 34207 21981
rect 33888 21944 33916 21975
rect 34974 21972 34980 21984
rect 35032 21972 35038 22024
rect 30708 21916 31340 21944
rect 31404 21916 33916 21944
rect 30708 21904 30714 21916
rect 11238 21836 11244 21888
rect 11296 21876 11302 21888
rect 12821 21879 12879 21885
rect 12821 21876 12833 21879
rect 11296 21848 12833 21876
rect 11296 21836 11302 21848
rect 12821 21845 12833 21848
rect 12867 21845 12879 21879
rect 12821 21839 12879 21845
rect 12989 21879 13047 21885
rect 12989 21845 13001 21879
rect 13035 21876 13047 21879
rect 13078 21876 13084 21888
rect 13035 21848 13084 21876
rect 13035 21845 13047 21848
rect 12989 21839 13047 21845
rect 13078 21836 13084 21848
rect 13136 21836 13142 21888
rect 15194 21836 15200 21888
rect 15252 21876 15258 21888
rect 16025 21879 16083 21885
rect 16025 21876 16037 21879
rect 15252 21848 16037 21876
rect 15252 21836 15258 21848
rect 16025 21845 16037 21848
rect 16071 21876 16083 21879
rect 16298 21876 16304 21888
rect 16071 21848 16304 21876
rect 16071 21845 16083 21848
rect 16025 21839 16083 21845
rect 16298 21836 16304 21848
rect 16356 21836 16362 21888
rect 16850 21836 16856 21888
rect 16908 21876 16914 21888
rect 17865 21879 17923 21885
rect 17865 21876 17877 21879
rect 16908 21848 17877 21876
rect 16908 21836 16914 21848
rect 17865 21845 17877 21848
rect 17911 21845 17923 21879
rect 17865 21839 17923 21845
rect 17954 21836 17960 21888
rect 18012 21876 18018 21888
rect 18525 21879 18583 21885
rect 18525 21876 18537 21879
rect 18012 21848 18537 21876
rect 18012 21836 18018 21848
rect 18525 21845 18537 21848
rect 18571 21845 18583 21879
rect 18690 21876 18696 21888
rect 18651 21848 18696 21876
rect 18525 21839 18583 21845
rect 18690 21836 18696 21848
rect 18748 21836 18754 21888
rect 21726 21836 21732 21888
rect 21784 21876 21790 21888
rect 21913 21879 21971 21885
rect 21913 21876 21925 21879
rect 21784 21848 21925 21876
rect 21784 21836 21790 21848
rect 21913 21845 21925 21848
rect 21959 21845 21971 21879
rect 23842 21876 23848 21888
rect 23755 21848 23848 21876
rect 21913 21839 21971 21845
rect 23842 21836 23848 21848
rect 23900 21876 23906 21888
rect 24578 21876 24584 21888
rect 23900 21848 24584 21876
rect 23900 21836 23906 21848
rect 24578 21836 24584 21848
rect 24636 21836 24642 21888
rect 25225 21879 25283 21885
rect 25225 21845 25237 21879
rect 25271 21876 25283 21879
rect 25314 21876 25320 21888
rect 25271 21848 25320 21876
rect 25271 21845 25283 21848
rect 25225 21839 25283 21845
rect 25314 21836 25320 21848
rect 25372 21836 25378 21888
rect 25774 21836 25780 21888
rect 25832 21836 25838 21888
rect 26329 21879 26387 21885
rect 26329 21845 26341 21879
rect 26375 21876 26387 21879
rect 31404 21876 31432 21916
rect 26375 21848 31432 21876
rect 32493 21879 32551 21885
rect 26375 21845 26387 21848
rect 26329 21839 26387 21845
rect 32493 21845 32505 21879
rect 32539 21876 32551 21879
rect 32766 21876 32772 21888
rect 32539 21848 32772 21876
rect 32539 21845 32551 21848
rect 32493 21839 32551 21845
rect 32766 21836 32772 21848
rect 32824 21836 32830 21888
rect 33689 21879 33747 21885
rect 33689 21845 33701 21879
rect 33735 21876 33747 21879
rect 33778 21876 33784 21888
rect 33735 21848 33784 21876
rect 33735 21845 33747 21848
rect 33689 21839 33747 21845
rect 33778 21836 33784 21848
rect 33836 21836 33842 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 7558 21632 7564 21684
rect 7616 21672 7622 21684
rect 7834 21672 7840 21684
rect 7892 21681 7898 21684
rect 7892 21675 7911 21681
rect 7616 21644 7840 21672
rect 7616 21632 7622 21644
rect 7834 21632 7840 21644
rect 7899 21672 7911 21675
rect 8481 21675 8539 21681
rect 8481 21672 8493 21675
rect 7899 21644 8493 21672
rect 7899 21641 7911 21644
rect 7892 21635 7911 21641
rect 8481 21641 8493 21644
rect 8527 21641 8539 21675
rect 8481 21635 8539 21641
rect 7892 21632 7898 21635
rect 12802 21632 12808 21684
rect 12860 21672 12866 21684
rect 12897 21675 12955 21681
rect 12897 21672 12909 21675
rect 12860 21644 12909 21672
rect 12860 21632 12866 21644
rect 12897 21641 12909 21644
rect 12943 21641 12955 21675
rect 15562 21672 15568 21684
rect 15523 21644 15568 21672
rect 12897 21635 12955 21641
rect 15562 21632 15568 21644
rect 15620 21632 15626 21684
rect 15654 21632 15660 21684
rect 15712 21672 15718 21684
rect 18598 21672 18604 21684
rect 15712 21644 18604 21672
rect 15712 21632 15718 21644
rect 18598 21632 18604 21644
rect 18656 21632 18662 21684
rect 18782 21672 18788 21684
rect 18743 21644 18788 21672
rect 18782 21632 18788 21644
rect 18840 21632 18846 21684
rect 19058 21632 19064 21684
rect 19116 21672 19122 21684
rect 22281 21675 22339 21681
rect 19116 21644 21956 21672
rect 19116 21632 19122 21644
rect 7374 21564 7380 21616
rect 7432 21604 7438 21616
rect 7653 21607 7711 21613
rect 7653 21604 7665 21607
rect 7432 21576 7665 21604
rect 7432 21564 7438 21576
rect 7653 21573 7665 21576
rect 7699 21573 7711 21607
rect 7653 21567 7711 21573
rect 11784 21607 11842 21613
rect 11784 21573 11796 21607
rect 11830 21604 11842 21607
rect 12342 21604 12348 21616
rect 11830 21576 12348 21604
rect 11830 21573 11842 21576
rect 11784 21567 11842 21573
rect 12342 21564 12348 21576
rect 12400 21564 12406 21616
rect 15105 21607 15163 21613
rect 15105 21573 15117 21607
rect 15151 21604 15163 21607
rect 15151 21576 16068 21604
rect 15151 21573 15163 21576
rect 15105 21567 15163 21573
rect 4433 21539 4491 21545
rect 4433 21505 4445 21539
rect 4479 21505 4491 21539
rect 5074 21536 5080 21548
rect 5035 21508 5080 21536
rect 4433 21499 4491 21505
rect 4448 21468 4476 21499
rect 5074 21496 5080 21508
rect 5132 21496 5138 21548
rect 6365 21539 6423 21545
rect 6365 21505 6377 21539
rect 6411 21536 6423 21539
rect 7006 21536 7012 21548
rect 6411 21508 7012 21536
rect 6411 21505 6423 21508
rect 6365 21499 6423 21505
rect 7006 21496 7012 21508
rect 7064 21496 7070 21548
rect 8662 21536 8668 21548
rect 8623 21508 8668 21536
rect 8662 21496 8668 21508
rect 8720 21496 8726 21548
rect 9214 21536 9220 21548
rect 9175 21508 9220 21536
rect 9214 21496 9220 21508
rect 9272 21496 9278 21548
rect 14918 21536 14924 21548
rect 14879 21508 14924 21536
rect 14918 21496 14924 21508
rect 14976 21496 14982 21548
rect 15746 21536 15752 21548
rect 15707 21508 15752 21536
rect 15746 21496 15752 21508
rect 15804 21496 15810 21548
rect 15838 21496 15844 21548
rect 15896 21536 15902 21548
rect 16040 21545 16068 21576
rect 16482 21564 16488 21616
rect 16540 21604 16546 21616
rect 16761 21607 16819 21613
rect 16761 21604 16773 21607
rect 16540 21576 16773 21604
rect 16540 21564 16546 21576
rect 16761 21573 16773 21576
rect 16807 21604 16819 21607
rect 19242 21604 19248 21616
rect 16807 21576 19248 21604
rect 16807 21573 16819 21576
rect 16761 21567 16819 21573
rect 19242 21564 19248 21576
rect 19300 21564 19306 21616
rect 21928 21613 21956 21644
rect 22281 21641 22293 21675
rect 22327 21672 22339 21675
rect 22646 21672 22652 21684
rect 22327 21644 22652 21672
rect 22327 21641 22339 21644
rect 22281 21635 22339 21641
rect 22646 21632 22652 21644
rect 22704 21632 22710 21684
rect 22830 21672 22836 21684
rect 22791 21644 22836 21672
rect 22830 21632 22836 21644
rect 22888 21632 22894 21684
rect 23106 21632 23112 21684
rect 23164 21672 23170 21684
rect 23164 21644 23244 21672
rect 23164 21632 23170 21644
rect 21913 21607 21971 21613
rect 21913 21573 21925 21607
rect 21959 21573 21971 21607
rect 21913 21567 21971 21573
rect 22129 21607 22187 21613
rect 22129 21573 22141 21607
rect 22175 21604 22187 21607
rect 22738 21604 22744 21616
rect 22175 21576 22744 21604
rect 22175 21573 22187 21576
rect 22129 21567 22187 21573
rect 22738 21564 22744 21576
rect 22796 21564 22802 21616
rect 23216 21604 23244 21644
rect 25038 21632 25044 21684
rect 25096 21672 25102 21684
rect 25317 21675 25375 21681
rect 25317 21672 25329 21675
rect 25096 21644 25329 21672
rect 25096 21632 25102 21644
rect 25317 21641 25329 21644
rect 25363 21641 25375 21675
rect 25317 21635 25375 21641
rect 27433 21675 27491 21681
rect 27433 21641 27445 21675
rect 27479 21672 27491 21675
rect 27706 21672 27712 21684
rect 27479 21644 27712 21672
rect 27479 21641 27491 21644
rect 27433 21635 27491 21641
rect 27706 21632 27712 21644
rect 27764 21632 27770 21684
rect 28258 21672 28264 21684
rect 27908 21644 28264 21672
rect 23658 21604 23664 21616
rect 23216 21576 23664 21604
rect 16025 21539 16083 21545
rect 15896 21508 15941 21536
rect 15896 21496 15902 21508
rect 16025 21505 16037 21539
rect 16071 21505 16083 21539
rect 16025 21499 16083 21505
rect 16117 21539 16175 21545
rect 16117 21505 16129 21539
rect 16163 21505 16175 21539
rect 16117 21499 16175 21505
rect 5718 21468 5724 21480
rect 4448 21440 5724 21468
rect 5718 21428 5724 21440
rect 5776 21428 5782 21480
rect 6454 21428 6460 21480
rect 6512 21468 6518 21480
rect 6641 21471 6699 21477
rect 6641 21468 6653 21471
rect 6512 21440 6653 21468
rect 6512 21428 6518 21440
rect 6641 21437 6653 21440
rect 6687 21437 6699 21471
rect 6641 21431 6699 21437
rect 10870 21428 10876 21480
rect 10928 21468 10934 21480
rect 11517 21471 11575 21477
rect 11517 21468 11529 21471
rect 10928 21440 11529 21468
rect 10928 21428 10934 21440
rect 11517 21437 11529 21440
rect 11563 21437 11575 21471
rect 11517 21431 11575 21437
rect 14737 21471 14795 21477
rect 14737 21437 14749 21471
rect 14783 21468 14795 21471
rect 15194 21468 15200 21480
rect 14783 21440 15200 21468
rect 14783 21437 14795 21440
rect 14737 21431 14795 21437
rect 15194 21428 15200 21440
rect 15252 21428 15258 21480
rect 16132 21468 16160 21499
rect 17310 21496 17316 21548
rect 17368 21536 17374 21548
rect 17405 21539 17463 21545
rect 17405 21536 17417 21539
rect 17368 21508 17417 21536
rect 17368 21496 17374 21508
rect 17405 21505 17417 21508
rect 17451 21505 17463 21539
rect 17405 21499 17463 21505
rect 17672 21539 17730 21545
rect 17672 21505 17684 21539
rect 17718 21536 17730 21539
rect 18414 21536 18420 21548
rect 17718 21508 18420 21536
rect 17718 21505 17730 21508
rect 17672 21499 17730 21505
rect 18414 21496 18420 21508
rect 18472 21496 18478 21548
rect 18690 21496 18696 21548
rect 18748 21536 18754 21548
rect 23216 21545 23244 21576
rect 23658 21564 23664 21576
rect 23716 21564 23722 21616
rect 27908 21604 27936 21644
rect 28258 21632 28264 21644
rect 28316 21632 28322 21684
rect 29914 21632 29920 21684
rect 29972 21672 29978 21684
rect 29972 21644 30052 21672
rect 29972 21632 29978 21644
rect 27448 21576 27936 21604
rect 28169 21607 28227 21613
rect 27448 21548 27476 21576
rect 28169 21573 28181 21607
rect 28215 21604 28227 21607
rect 28276 21604 28304 21632
rect 28215 21576 28304 21604
rect 28215 21573 28227 21576
rect 28169 21567 28227 21573
rect 28442 21564 28448 21616
rect 28500 21604 28506 21616
rect 29546 21604 29552 21616
rect 28500 21576 29552 21604
rect 28500 21564 28506 21576
rect 29546 21564 29552 21576
rect 29604 21564 29610 21616
rect 19429 21539 19487 21545
rect 19429 21536 19441 21539
rect 18748 21508 19441 21536
rect 18748 21496 18754 21508
rect 19429 21505 19441 21508
rect 19475 21505 19487 21539
rect 23109 21539 23167 21545
rect 23109 21536 23121 21539
rect 19429 21499 19487 21505
rect 23032 21508 23121 21536
rect 16758 21468 16764 21480
rect 16132 21440 16764 21468
rect 9490 21400 9496 21412
rect 7852 21372 9496 21400
rect 4249 21335 4307 21341
rect 4249 21301 4261 21335
rect 4295 21332 4307 21335
rect 4614 21332 4620 21344
rect 4295 21304 4620 21332
rect 4295 21301 4307 21304
rect 4249 21295 4307 21301
rect 4614 21292 4620 21304
rect 4672 21292 4678 21344
rect 4890 21332 4896 21344
rect 4851 21304 4896 21332
rect 4890 21292 4896 21304
rect 4948 21292 4954 21344
rect 7852 21341 7880 21372
rect 9490 21360 9496 21372
rect 9548 21360 9554 21412
rect 15562 21360 15568 21412
rect 15620 21400 15626 21412
rect 16132 21400 16160 21440
rect 16758 21428 16764 21440
rect 16816 21428 16822 21480
rect 16945 21471 17003 21477
rect 16945 21437 16957 21471
rect 16991 21468 17003 21471
rect 17126 21468 17132 21480
rect 16991 21440 17132 21468
rect 16991 21437 17003 21440
rect 16945 21431 17003 21437
rect 17126 21428 17132 21440
rect 17184 21428 17190 21480
rect 19705 21471 19763 21477
rect 19705 21437 19717 21471
rect 19751 21468 19763 21471
rect 20898 21468 20904 21480
rect 19751 21440 20904 21468
rect 19751 21437 19763 21440
rect 19705 21431 19763 21437
rect 20898 21428 20904 21440
rect 20956 21428 20962 21480
rect 15620 21372 16160 21400
rect 23032 21400 23060 21508
rect 23109 21505 23121 21508
rect 23155 21505 23167 21539
rect 23109 21499 23167 21505
rect 23201 21539 23259 21545
rect 23201 21505 23213 21539
rect 23247 21505 23259 21539
rect 23201 21499 23259 21505
rect 23293 21539 23351 21545
rect 23293 21505 23305 21539
rect 23339 21505 23351 21539
rect 23293 21499 23351 21505
rect 23308 21468 23336 21499
rect 23382 21496 23388 21548
rect 23440 21536 23446 21548
rect 23477 21539 23535 21545
rect 23477 21536 23489 21539
rect 23440 21508 23489 21536
rect 23440 21496 23446 21508
rect 23477 21505 23489 21508
rect 23523 21505 23535 21539
rect 24026 21536 24032 21548
rect 23987 21508 24032 21536
rect 23477 21499 23535 21505
rect 24026 21496 24032 21508
rect 24084 21496 24090 21548
rect 27065 21539 27123 21545
rect 27065 21505 27077 21539
rect 27111 21536 27123 21539
rect 27154 21536 27160 21548
rect 27111 21508 27160 21536
rect 27111 21505 27123 21508
rect 27065 21499 27123 21505
rect 27154 21496 27160 21508
rect 27212 21496 27218 21548
rect 27249 21539 27307 21545
rect 27249 21505 27261 21539
rect 27295 21505 27307 21539
rect 27249 21499 27307 21505
rect 23658 21468 23664 21480
rect 23308 21440 23664 21468
rect 23658 21428 23664 21440
rect 23716 21428 23722 21480
rect 27264 21468 27292 21499
rect 27430 21496 27436 21548
rect 27488 21496 27494 21548
rect 27890 21536 27896 21548
rect 27851 21508 27896 21536
rect 27890 21496 27896 21508
rect 27948 21496 27954 21548
rect 27986 21539 28044 21545
rect 27986 21505 27998 21539
rect 28032 21505 28044 21539
rect 27986 21499 28044 21505
rect 28261 21539 28319 21545
rect 28261 21505 28273 21539
rect 28307 21505 28319 21539
rect 28261 21499 28319 21505
rect 27264 21440 27614 21468
rect 24578 21400 24584 21412
rect 23032 21372 24584 21400
rect 15620 21360 15626 21372
rect 24578 21360 24584 21372
rect 24636 21360 24642 21412
rect 27586 21400 27614 21440
rect 27998 21400 28026 21499
rect 28074 21400 28080 21412
rect 27586 21372 28080 21400
rect 28074 21360 28080 21372
rect 28132 21360 28138 21412
rect 28276 21400 28304 21499
rect 28350 21496 28356 21548
rect 28408 21545 28414 21548
rect 28408 21536 28416 21545
rect 28994 21536 29000 21548
rect 28408 21508 28453 21536
rect 28955 21508 29000 21536
rect 28408 21499 28416 21508
rect 28408 21496 28414 21499
rect 28994 21496 29000 21508
rect 29052 21496 29058 21548
rect 29181 21539 29239 21545
rect 29181 21505 29193 21539
rect 29227 21536 29239 21539
rect 29270 21536 29276 21548
rect 29227 21508 29276 21536
rect 29227 21505 29239 21508
rect 29181 21499 29239 21505
rect 29270 21496 29276 21508
rect 29328 21496 29334 21548
rect 29730 21496 29736 21548
rect 29788 21536 29794 21548
rect 30024 21545 30052 21644
rect 30098 21632 30104 21684
rect 30156 21672 30162 21684
rect 31021 21675 31079 21681
rect 30156 21644 30420 21672
rect 30156 21632 30162 21644
rect 30208 21613 30236 21644
rect 30193 21607 30251 21613
rect 30193 21573 30205 21607
rect 30239 21573 30251 21607
rect 30392 21604 30420 21644
rect 31021 21641 31033 21675
rect 31067 21672 31079 21675
rect 31570 21672 31576 21684
rect 31067 21644 31576 21672
rect 31067 21641 31079 21644
rect 31021 21635 31079 21641
rect 31570 21632 31576 21644
rect 31628 21632 31634 21684
rect 32674 21672 32680 21684
rect 32635 21644 32680 21672
rect 32674 21632 32680 21644
rect 32732 21632 32738 21684
rect 34974 21672 34980 21684
rect 34935 21644 34980 21672
rect 34974 21632 34980 21644
rect 35032 21632 35038 21684
rect 32309 21607 32367 21613
rect 30392 21576 31156 21604
rect 30193 21567 30251 21573
rect 29825 21539 29883 21545
rect 29825 21536 29837 21539
rect 29788 21508 29837 21536
rect 29788 21496 29794 21508
rect 29825 21505 29837 21508
rect 29871 21505 29883 21539
rect 29825 21499 29883 21505
rect 29973 21539 30052 21545
rect 29973 21505 29985 21539
rect 30019 21508 30052 21539
rect 30019 21505 30031 21508
rect 29973 21499 30031 21505
rect 30098 21496 30104 21548
rect 30156 21536 30162 21548
rect 30331 21539 30389 21545
rect 30156 21508 30201 21536
rect 30156 21496 30162 21508
rect 30331 21505 30343 21539
rect 30377 21536 30389 21539
rect 30466 21536 30472 21548
rect 30377 21508 30472 21536
rect 30377 21505 30389 21508
rect 30331 21499 30389 21505
rect 30466 21496 30472 21508
rect 30524 21496 30530 21548
rect 30926 21536 30932 21548
rect 30887 21508 30932 21536
rect 30926 21496 30932 21508
rect 30984 21496 30990 21548
rect 31128 21545 31156 21576
rect 32309 21573 32321 21607
rect 32355 21604 32367 21607
rect 33502 21604 33508 21616
rect 32355 21576 33508 21604
rect 32355 21573 32367 21576
rect 32309 21567 32367 21573
rect 33502 21564 33508 21576
rect 33560 21564 33566 21616
rect 33864 21607 33922 21613
rect 33864 21573 33876 21607
rect 33910 21604 33922 21607
rect 33962 21604 33968 21616
rect 33910 21576 33968 21604
rect 33910 21573 33922 21576
rect 33864 21567 33922 21573
rect 33962 21564 33968 21576
rect 34020 21564 34026 21616
rect 31113 21539 31171 21545
rect 31113 21505 31125 21539
rect 31159 21536 31171 21539
rect 31938 21536 31944 21548
rect 31159 21508 31944 21536
rect 31159 21505 31171 21508
rect 31113 21499 31171 21505
rect 31938 21496 31944 21508
rect 31996 21496 32002 21548
rect 32493 21539 32551 21545
rect 32493 21505 32505 21539
rect 32539 21536 32551 21539
rect 32766 21536 32772 21548
rect 32539 21508 32772 21536
rect 32539 21505 32551 21508
rect 32493 21499 32551 21505
rect 32766 21496 32772 21508
rect 32824 21496 32830 21548
rect 29365 21471 29423 21477
rect 29365 21437 29377 21471
rect 29411 21468 29423 21471
rect 31386 21468 31392 21480
rect 29411 21440 31392 21468
rect 29411 21437 29423 21440
rect 29365 21431 29423 21437
rect 31386 21428 31392 21440
rect 31444 21428 31450 21480
rect 33594 21468 33600 21480
rect 33555 21440 33600 21468
rect 33594 21428 33600 21440
rect 33652 21428 33658 21480
rect 31202 21400 31208 21412
rect 28276 21372 31208 21400
rect 31202 21360 31208 21372
rect 31260 21360 31266 21412
rect 7837 21335 7895 21341
rect 7837 21301 7849 21335
rect 7883 21301 7895 21335
rect 7837 21295 7895 21301
rect 8021 21335 8079 21341
rect 8021 21301 8033 21335
rect 8067 21332 8079 21335
rect 8294 21332 8300 21344
rect 8067 21304 8300 21332
rect 8067 21301 8079 21304
rect 8021 21295 8079 21301
rect 8294 21292 8300 21304
rect 8352 21292 8358 21344
rect 8938 21292 8944 21344
rect 8996 21332 9002 21344
rect 10505 21335 10563 21341
rect 10505 21332 10517 21335
rect 8996 21304 10517 21332
rect 8996 21292 9002 21304
rect 10505 21301 10517 21304
rect 10551 21301 10563 21335
rect 10505 21295 10563 21301
rect 22094 21292 22100 21344
rect 22152 21332 22158 21344
rect 22152 21304 22197 21332
rect 22152 21292 22158 21304
rect 24394 21292 24400 21344
rect 24452 21332 24458 21344
rect 25590 21332 25596 21344
rect 24452 21304 25596 21332
rect 24452 21292 24458 21304
rect 25590 21292 25596 21304
rect 25648 21332 25654 21344
rect 27062 21332 27068 21344
rect 25648 21304 27068 21332
rect 25648 21292 25654 21304
rect 27062 21292 27068 21304
rect 27120 21292 27126 21344
rect 28258 21292 28264 21344
rect 28316 21332 28322 21344
rect 28537 21335 28595 21341
rect 28537 21332 28549 21335
rect 28316 21304 28549 21332
rect 28316 21292 28322 21304
rect 28537 21301 28549 21304
rect 28583 21301 28595 21335
rect 30466 21332 30472 21344
rect 30427 21304 30472 21332
rect 28537 21295 28595 21301
rect 30466 21292 30472 21304
rect 30524 21292 30530 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 6270 21128 6276 21140
rect 6231 21100 6276 21128
rect 6270 21088 6276 21100
rect 6328 21088 6334 21140
rect 7561 21131 7619 21137
rect 7561 21097 7573 21131
rect 7607 21097 7619 21131
rect 7561 21091 7619 21097
rect 7745 21131 7803 21137
rect 7745 21097 7757 21131
rect 7791 21128 7803 21131
rect 9582 21128 9588 21140
rect 7791 21100 9588 21128
rect 7791 21097 7803 21100
rect 7745 21091 7803 21097
rect 3786 20924 3792 20936
rect 3747 20896 3792 20924
rect 3786 20884 3792 20896
rect 3844 20884 3850 20936
rect 4056 20927 4114 20933
rect 4056 20893 4068 20927
rect 4102 20924 4114 20927
rect 4890 20924 4896 20936
rect 4102 20896 4896 20924
rect 4102 20893 4114 20896
rect 4056 20887 4114 20893
rect 4890 20884 4896 20896
rect 4948 20884 4954 20936
rect 6457 20927 6515 20933
rect 6457 20893 6469 20927
rect 6503 20924 6515 20927
rect 6914 20924 6920 20936
rect 6503 20896 6920 20924
rect 6503 20893 6515 20896
rect 6457 20887 6515 20893
rect 6914 20884 6920 20896
rect 6972 20884 6978 20936
rect 7374 20856 7380 20868
rect 7335 20828 7380 20856
rect 7374 20816 7380 20828
rect 7432 20816 7438 20868
rect 7576 20856 7604 21091
rect 9582 21088 9588 21100
rect 9640 21088 9646 21140
rect 11330 21128 11336 21140
rect 11291 21100 11336 21128
rect 11330 21088 11336 21100
rect 11388 21088 11394 21140
rect 12710 21088 12716 21140
rect 12768 21128 12774 21140
rect 12805 21131 12863 21137
rect 12805 21128 12817 21131
rect 12768 21100 12817 21128
rect 12768 21088 12774 21100
rect 12805 21097 12817 21100
rect 12851 21097 12863 21131
rect 16206 21128 16212 21140
rect 16167 21100 16212 21128
rect 12805 21091 12863 21097
rect 16206 21088 16212 21100
rect 16264 21088 16270 21140
rect 18414 21128 18420 21140
rect 18375 21100 18420 21128
rect 18414 21088 18420 21100
rect 18472 21088 18478 21140
rect 22278 21088 22284 21140
rect 22336 21128 22342 21140
rect 22649 21131 22707 21137
rect 22649 21128 22661 21131
rect 22336 21100 22661 21128
rect 22336 21088 22342 21100
rect 22649 21097 22661 21100
rect 22695 21097 22707 21131
rect 22649 21091 22707 21097
rect 23477 21131 23535 21137
rect 23477 21097 23489 21131
rect 23523 21128 23535 21131
rect 23658 21128 23664 21140
rect 23523 21100 23664 21128
rect 23523 21097 23535 21100
rect 23477 21091 23535 21097
rect 23658 21088 23664 21100
rect 23716 21088 23722 21140
rect 25130 21128 25136 21140
rect 23768 21100 25136 21128
rect 21266 21060 21272 21072
rect 21008 21032 21272 21060
rect 8938 20992 8944 21004
rect 8899 20964 8944 20992
rect 8938 20952 8944 20964
rect 8996 20952 9002 21004
rect 14090 20992 14096 21004
rect 14051 20964 14096 20992
rect 14090 20952 14096 20964
rect 14148 20952 14154 21004
rect 15378 20952 15384 21004
rect 15436 20992 15442 21004
rect 15838 20992 15844 21004
rect 15436 20964 15844 20992
rect 15436 20952 15442 20964
rect 15838 20952 15844 20964
rect 15896 20992 15902 21004
rect 21008 21001 21036 21032
rect 21266 21020 21272 21032
rect 21324 21020 21330 21072
rect 20993 20995 21051 21001
rect 15896 20964 16528 20992
rect 15896 20952 15902 20964
rect 8389 20927 8447 20933
rect 8389 20893 8401 20927
rect 8435 20924 8447 20927
rect 8478 20924 8484 20936
rect 8435 20896 8484 20924
rect 8435 20893 8447 20896
rect 8389 20887 8447 20893
rect 8478 20884 8484 20896
rect 8536 20884 8542 20936
rect 11517 20927 11575 20933
rect 11517 20893 11529 20927
rect 11563 20924 11575 20927
rect 11882 20924 11888 20936
rect 11563 20896 11888 20924
rect 11563 20893 11575 20896
rect 11517 20887 11575 20893
rect 11882 20884 11888 20896
rect 11940 20884 11946 20936
rect 12713 20927 12771 20933
rect 12713 20893 12725 20927
rect 12759 20924 12771 20927
rect 12894 20924 12900 20936
rect 12759 20896 12900 20924
rect 12759 20893 12771 20896
rect 12713 20887 12771 20893
rect 12894 20884 12900 20896
rect 12952 20884 12958 20936
rect 13814 20884 13820 20936
rect 13872 20884 13878 20936
rect 16500 20933 16528 20964
rect 20993 20961 21005 20995
rect 21039 20961 21051 20995
rect 20993 20955 21051 20961
rect 16393 20927 16451 20933
rect 16393 20893 16405 20927
rect 16439 20893 16451 20927
rect 16393 20887 16451 20893
rect 16485 20927 16543 20933
rect 16485 20893 16497 20927
rect 16531 20893 16543 20927
rect 16666 20924 16672 20936
rect 16627 20896 16672 20924
rect 16485 20887 16543 20893
rect 9208 20859 9266 20865
rect 7576 20828 9168 20856
rect 4798 20748 4804 20800
rect 4856 20788 4862 20800
rect 5169 20791 5227 20797
rect 5169 20788 5181 20791
rect 4856 20760 5181 20788
rect 4856 20748 4862 20760
rect 5169 20757 5181 20760
rect 5215 20757 5227 20791
rect 5169 20751 5227 20757
rect 7558 20748 7564 20800
rect 7616 20797 7622 20800
rect 7616 20791 7635 20797
rect 7623 20757 7635 20791
rect 7616 20751 7635 20757
rect 8205 20791 8263 20797
rect 8205 20757 8217 20791
rect 8251 20788 8263 20791
rect 9030 20788 9036 20800
rect 8251 20760 9036 20788
rect 8251 20757 8263 20760
rect 8205 20751 8263 20757
rect 7616 20748 7622 20751
rect 9030 20748 9036 20760
rect 9088 20748 9094 20800
rect 9140 20788 9168 20828
rect 9208 20825 9220 20859
rect 9254 20856 9266 20859
rect 10410 20856 10416 20868
rect 9254 20828 10416 20856
rect 9254 20825 9266 20828
rect 9208 20819 9266 20825
rect 10410 20816 10416 20828
rect 10468 20816 10474 20868
rect 13832 20856 13860 20884
rect 14090 20856 14096 20868
rect 13832 20828 14096 20856
rect 14090 20816 14096 20828
rect 14148 20816 14154 20868
rect 14360 20859 14418 20865
rect 14360 20825 14372 20859
rect 14406 20856 14418 20859
rect 14734 20856 14740 20868
rect 14406 20828 14740 20856
rect 14406 20825 14418 20828
rect 14360 20819 14418 20825
rect 14734 20816 14740 20828
rect 14792 20816 14798 20868
rect 16408 20856 16436 20887
rect 16666 20884 16672 20896
rect 16724 20884 16730 20936
rect 16758 20884 16764 20936
rect 16816 20924 16822 20936
rect 17770 20924 17776 20936
rect 16816 20896 16988 20924
rect 17731 20896 17776 20924
rect 16816 20884 16822 20896
rect 16574 20856 16580 20868
rect 16408 20828 16580 20856
rect 16574 20816 16580 20828
rect 16632 20856 16638 20868
rect 16960 20856 16988 20896
rect 17770 20884 17776 20896
rect 17828 20884 17834 20936
rect 19245 20927 19303 20933
rect 19245 20893 19257 20927
rect 19291 20924 19303 20927
rect 19426 20924 19432 20936
rect 19291 20896 19432 20924
rect 19291 20893 19303 20896
rect 19245 20887 19303 20893
rect 19426 20884 19432 20896
rect 19484 20884 19490 20936
rect 19521 20927 19579 20933
rect 19521 20893 19533 20927
rect 19567 20893 19579 20927
rect 19521 20887 19579 20893
rect 21269 20927 21327 20933
rect 21269 20893 21281 20927
rect 21315 20924 21327 20927
rect 22281 20927 22339 20933
rect 22281 20924 22293 20927
rect 21315 20896 22293 20924
rect 21315 20893 21327 20896
rect 21269 20887 21327 20893
rect 22281 20893 22293 20896
rect 22327 20924 22339 20927
rect 23109 20927 23167 20933
rect 23109 20924 23121 20927
rect 22327 20896 23121 20924
rect 22327 20893 22339 20896
rect 22281 20887 22339 20893
rect 23109 20893 23121 20896
rect 23155 20924 23167 20927
rect 23768 20924 23796 21100
rect 25130 21088 25136 21100
rect 25188 21088 25194 21140
rect 25314 21088 25320 21140
rect 25372 21128 25378 21140
rect 29917 21131 29975 21137
rect 25372 21100 28028 21128
rect 25372 21088 25378 21100
rect 24670 21020 24676 21072
rect 24728 21060 24734 21072
rect 26513 21063 26571 21069
rect 26513 21060 26525 21063
rect 24728 21032 26525 21060
rect 24728 21020 24734 21032
rect 26513 21029 26525 21032
rect 26559 21060 26571 21063
rect 26970 21060 26976 21072
rect 26559 21032 26976 21060
rect 26559 21029 26571 21032
rect 26513 21023 26571 21029
rect 26970 21020 26976 21032
rect 27028 21020 27034 21072
rect 27249 21063 27307 21069
rect 27249 21029 27261 21063
rect 27295 21060 27307 21063
rect 27706 21060 27712 21072
rect 27295 21032 27712 21060
rect 27295 21029 27307 21032
rect 27249 21023 27307 21029
rect 27706 21020 27712 21032
rect 27764 21020 27770 21072
rect 28000 21060 28028 21100
rect 29917 21097 29929 21131
rect 29963 21128 29975 21131
rect 30282 21128 30288 21140
rect 29963 21100 30288 21128
rect 29963 21097 29975 21100
rect 29917 21091 29975 21097
rect 30282 21088 30288 21100
rect 30340 21088 30346 21140
rect 31754 21128 31760 21140
rect 30392 21100 31760 21128
rect 30392 21060 30420 21100
rect 31754 21088 31760 21100
rect 31812 21088 31818 21140
rect 31938 21128 31944 21140
rect 31899 21100 31944 21128
rect 31938 21088 31944 21100
rect 31996 21088 32002 21140
rect 33965 21131 34023 21137
rect 33965 21097 33977 21131
rect 34011 21128 34023 21131
rect 34146 21128 34152 21140
rect 34011 21100 34152 21128
rect 34011 21097 34023 21100
rect 33965 21091 34023 21097
rect 34146 21088 34152 21100
rect 34204 21088 34210 21140
rect 28000 21032 30420 21060
rect 25130 20952 25136 21004
rect 25188 20992 25194 21004
rect 25188 20964 27844 20992
rect 25188 20952 25194 20964
rect 24394 20924 24400 20936
rect 23155 20896 23796 20924
rect 24228 20896 24400 20924
rect 23155 20893 23167 20896
rect 23109 20887 23167 20893
rect 18230 20856 18236 20868
rect 16632 20828 16896 20856
rect 16960 20828 18236 20856
rect 16632 20816 16638 20828
rect 10321 20791 10379 20797
rect 10321 20788 10333 20791
rect 9140 20760 10333 20788
rect 10321 20757 10333 20760
rect 10367 20757 10379 20791
rect 10321 20751 10379 20757
rect 13814 20748 13820 20800
rect 13872 20788 13878 20800
rect 15473 20791 15531 20797
rect 15473 20788 15485 20791
rect 13872 20760 15485 20788
rect 13872 20748 13878 20760
rect 15473 20757 15485 20760
rect 15519 20757 15531 20791
rect 16868 20788 16896 20828
rect 18230 20816 18236 20828
rect 18288 20816 18294 20868
rect 19536 20856 19564 20887
rect 19306 20828 19564 20856
rect 22465 20859 22523 20865
rect 19306 20800 19334 20828
rect 22465 20825 22477 20859
rect 22511 20856 22523 20859
rect 22646 20856 22652 20868
rect 22511 20828 22652 20856
rect 22511 20825 22523 20828
rect 22465 20819 22523 20825
rect 22646 20816 22652 20828
rect 22704 20816 22710 20868
rect 23290 20856 23296 20868
rect 23251 20828 23296 20856
rect 23290 20816 23296 20828
rect 23348 20816 23354 20868
rect 17218 20788 17224 20800
rect 16868 20760 17224 20788
rect 15473 20751 15531 20757
rect 17218 20748 17224 20760
rect 17276 20748 17282 20800
rect 18322 20748 18328 20800
rect 18380 20788 18386 20800
rect 18690 20788 18696 20800
rect 18380 20760 18696 20788
rect 18380 20748 18386 20760
rect 18690 20748 18696 20760
rect 18748 20748 18754 20800
rect 19242 20748 19248 20800
rect 19300 20760 19334 20800
rect 19300 20748 19306 20760
rect 19426 20748 19432 20800
rect 19484 20788 19490 20800
rect 24228 20788 24256 20896
rect 24394 20884 24400 20896
rect 24452 20884 24458 20936
rect 24490 20927 24548 20933
rect 24490 20893 24502 20927
rect 24536 20893 24548 20927
rect 24490 20887 24548 20893
rect 24302 20816 24308 20868
rect 24360 20856 24366 20868
rect 24505 20856 24533 20887
rect 24578 20884 24584 20936
rect 24636 20924 24642 20936
rect 24765 20927 24823 20933
rect 24765 20924 24777 20927
rect 24636 20896 24777 20924
rect 24636 20884 24642 20896
rect 24765 20893 24777 20896
rect 24811 20893 24823 20927
rect 24765 20887 24823 20893
rect 24903 20927 24961 20933
rect 24903 20893 24915 20927
rect 24949 20924 24961 20927
rect 26510 20924 26516 20936
rect 24949 20896 26516 20924
rect 24949 20893 24961 20896
rect 24903 20887 24961 20893
rect 26510 20884 26516 20896
rect 26568 20884 26574 20936
rect 27816 20933 27844 20964
rect 28166 20952 28172 21004
rect 28224 20992 28230 21004
rect 28224 20964 29776 20992
rect 28224 20952 28230 20964
rect 27801 20927 27859 20933
rect 27801 20893 27813 20927
rect 27847 20924 27859 20927
rect 28994 20924 29000 20936
rect 27847 20896 29000 20924
rect 27847 20893 27859 20896
rect 27801 20887 27859 20893
rect 28994 20884 29000 20896
rect 29052 20924 29058 20936
rect 29748 20933 29776 20964
rect 29822 20952 29828 21004
rect 29880 20992 29886 21004
rect 29880 20964 30696 20992
rect 29880 20952 29886 20964
rect 29549 20927 29607 20933
rect 29549 20924 29561 20927
rect 29052 20896 29561 20924
rect 29052 20884 29058 20896
rect 29549 20893 29561 20896
rect 29595 20893 29607 20927
rect 29549 20887 29607 20893
rect 29733 20927 29791 20933
rect 29733 20893 29745 20927
rect 29779 20893 29791 20927
rect 30558 20924 30564 20936
rect 30519 20896 30564 20924
rect 29733 20887 29791 20893
rect 30558 20884 30564 20896
rect 30616 20884 30622 20936
rect 30668 20924 30696 20964
rect 30817 20927 30875 20933
rect 30817 20924 30829 20927
rect 30668 20896 30829 20924
rect 30817 20893 30829 20896
rect 30863 20893 30875 20927
rect 30817 20887 30875 20893
rect 24670 20856 24676 20868
rect 24360 20828 24533 20856
rect 24631 20828 24676 20856
rect 24360 20816 24366 20828
rect 24670 20816 24676 20828
rect 24728 20816 24734 20868
rect 25593 20859 25651 20865
rect 25593 20825 25605 20859
rect 25639 20856 25651 20859
rect 25774 20856 25780 20868
rect 25639 20828 25780 20856
rect 25639 20825 25651 20828
rect 25593 20819 25651 20825
rect 25774 20816 25780 20828
rect 25832 20856 25838 20868
rect 26329 20859 26387 20865
rect 26329 20856 26341 20859
rect 25832 20828 26341 20856
rect 25832 20816 25838 20828
rect 26329 20825 26341 20828
rect 26375 20825 26387 20859
rect 26329 20819 26387 20825
rect 27062 20816 27068 20868
rect 27120 20856 27126 20868
rect 27985 20859 28043 20865
rect 27985 20856 27997 20859
rect 27120 20828 27165 20856
rect 27244 20828 27997 20856
rect 27120 20816 27126 20828
rect 19484 20760 24256 20788
rect 19484 20748 19490 20760
rect 24578 20748 24584 20800
rect 24636 20788 24642 20800
rect 25041 20791 25099 20797
rect 25041 20788 25053 20791
rect 24636 20760 25053 20788
rect 24636 20748 24642 20760
rect 25041 20757 25053 20760
rect 25087 20757 25099 20791
rect 25682 20788 25688 20800
rect 25643 20760 25688 20788
rect 25041 20751 25099 20757
rect 25682 20748 25688 20760
rect 25740 20748 25746 20800
rect 26602 20748 26608 20800
rect 26660 20788 26666 20800
rect 27244 20788 27272 20828
rect 27985 20825 27997 20828
rect 28031 20825 28043 20859
rect 27985 20819 28043 20825
rect 28074 20816 28080 20868
rect 28132 20856 28138 20868
rect 30098 20856 30104 20868
rect 28132 20828 30104 20856
rect 28132 20816 28138 20828
rect 30098 20816 30104 20828
rect 30156 20816 30162 20868
rect 33502 20816 33508 20868
rect 33560 20856 33566 20868
rect 33597 20859 33655 20865
rect 33597 20856 33609 20859
rect 33560 20828 33609 20856
rect 33560 20816 33566 20828
rect 33597 20825 33609 20828
rect 33643 20825 33655 20859
rect 33778 20856 33784 20868
rect 33739 20828 33784 20856
rect 33597 20819 33655 20825
rect 33778 20816 33784 20828
rect 33836 20816 33842 20868
rect 26660 20760 27272 20788
rect 28169 20791 28227 20797
rect 26660 20748 26666 20760
rect 28169 20757 28181 20791
rect 28215 20788 28227 20791
rect 28442 20788 28448 20800
rect 28215 20760 28448 20788
rect 28215 20757 28227 20760
rect 28169 20751 28227 20757
rect 28442 20748 28448 20760
rect 28500 20748 28506 20800
rect 28718 20748 28724 20800
rect 28776 20788 28782 20800
rect 29822 20788 29828 20800
rect 28776 20760 29828 20788
rect 28776 20748 28782 20760
rect 29822 20748 29828 20760
rect 29880 20748 29886 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 5534 20544 5540 20596
rect 5592 20593 5598 20596
rect 5592 20587 5611 20593
rect 5599 20553 5611 20587
rect 5718 20584 5724 20596
rect 5679 20556 5724 20584
rect 5592 20547 5611 20553
rect 5592 20544 5598 20547
rect 5718 20544 5724 20556
rect 5776 20544 5782 20596
rect 6565 20587 6623 20593
rect 6565 20584 6577 20587
rect 5828 20556 6577 20584
rect 3780 20519 3838 20525
rect 3780 20485 3792 20519
rect 3826 20516 3838 20519
rect 4614 20516 4620 20528
rect 3826 20488 4620 20516
rect 3826 20485 3838 20488
rect 3780 20479 3838 20485
rect 4614 20476 4620 20488
rect 4672 20476 4678 20528
rect 5353 20519 5411 20525
rect 5353 20485 5365 20519
rect 5399 20516 5411 20519
rect 5442 20516 5448 20528
rect 5399 20488 5448 20516
rect 5399 20485 5411 20488
rect 5353 20479 5411 20485
rect 5442 20476 5448 20488
rect 5500 20476 5506 20528
rect 5552 20516 5580 20544
rect 5828 20516 5856 20556
rect 6565 20553 6577 20556
rect 6611 20553 6623 20587
rect 6565 20547 6623 20553
rect 6733 20587 6791 20593
rect 6733 20553 6745 20587
rect 6779 20553 6791 20587
rect 10410 20584 10416 20596
rect 10371 20556 10416 20584
rect 6733 20547 6791 20553
rect 5552 20488 5856 20516
rect 5902 20476 5908 20528
rect 5960 20516 5966 20528
rect 6365 20519 6423 20525
rect 6365 20516 6377 20519
rect 5960 20488 6377 20516
rect 5960 20476 5966 20488
rect 6365 20485 6377 20488
rect 6411 20516 6423 20519
rect 6454 20516 6460 20528
rect 6411 20488 6460 20516
rect 6411 20485 6423 20488
rect 6365 20479 6423 20485
rect 6454 20476 6460 20488
rect 6512 20476 6518 20528
rect 3053 20451 3111 20457
rect 3053 20417 3065 20451
rect 3099 20448 3111 20451
rect 6748 20448 6776 20547
rect 10410 20544 10416 20556
rect 10468 20544 10474 20596
rect 11701 20587 11759 20593
rect 11701 20553 11713 20587
rect 11747 20584 11759 20587
rect 12894 20584 12900 20596
rect 11747 20556 12900 20584
rect 11747 20553 11759 20556
rect 11701 20547 11759 20553
rect 12894 20544 12900 20556
rect 12952 20544 12958 20596
rect 13906 20544 13912 20596
rect 13964 20584 13970 20596
rect 14366 20584 14372 20596
rect 13964 20556 14372 20584
rect 13964 20544 13970 20556
rect 14366 20544 14372 20556
rect 14424 20544 14430 20596
rect 14734 20584 14740 20596
rect 14695 20556 14740 20584
rect 14734 20544 14740 20556
rect 14792 20544 14798 20596
rect 15286 20544 15292 20596
rect 15344 20584 15350 20596
rect 15654 20584 15660 20596
rect 15344 20556 15660 20584
rect 15344 20544 15350 20556
rect 15654 20544 15660 20556
rect 15712 20544 15718 20596
rect 17681 20587 17739 20593
rect 15764 20556 16988 20584
rect 7374 20516 7380 20528
rect 7335 20488 7380 20516
rect 7374 20476 7380 20488
rect 7432 20476 7438 20528
rect 7558 20476 7564 20528
rect 7616 20525 7622 20528
rect 7616 20519 7635 20525
rect 7623 20485 7635 20519
rect 8938 20516 8944 20528
rect 7616 20479 7635 20485
rect 8588 20488 8944 20516
rect 7616 20476 7622 20479
rect 8588 20457 8616 20488
rect 8938 20476 8944 20488
rect 8996 20476 9002 20528
rect 14093 20519 14151 20525
rect 14093 20485 14105 20519
rect 14139 20516 14151 20519
rect 15764 20516 15792 20556
rect 16850 20516 16856 20528
rect 14139 20488 15792 20516
rect 15856 20488 16856 20516
rect 14139 20485 14151 20488
rect 14093 20479 14151 20485
rect 3099 20420 6776 20448
rect 8573 20451 8631 20457
rect 3099 20417 3111 20420
rect 3053 20411 3111 20417
rect 8573 20417 8585 20451
rect 8619 20417 8631 20451
rect 8573 20411 8631 20417
rect 8662 20408 8668 20460
rect 8720 20448 8726 20460
rect 8829 20451 8887 20457
rect 8829 20448 8841 20451
rect 8720 20420 8841 20448
rect 8720 20408 8726 20420
rect 8829 20417 8841 20420
rect 8875 20417 8887 20451
rect 8829 20411 8887 20417
rect 9582 20408 9588 20460
rect 9640 20448 9646 20460
rect 10597 20451 10655 20457
rect 10597 20448 10609 20451
rect 9640 20420 10609 20448
rect 9640 20408 9646 20420
rect 10597 20417 10609 20420
rect 10643 20417 10655 20451
rect 11514 20448 11520 20460
rect 11475 20420 11520 20448
rect 10597 20411 10655 20417
rect 11514 20408 11520 20420
rect 11572 20408 11578 20460
rect 13357 20451 13415 20457
rect 13357 20417 13369 20451
rect 13403 20448 13415 20451
rect 13814 20448 13820 20460
rect 13403 20420 13820 20448
rect 13403 20417 13415 20420
rect 13357 20411 13415 20417
rect 13814 20408 13820 20420
rect 13872 20408 13878 20460
rect 14642 20408 14648 20460
rect 14700 20448 14706 20460
rect 14918 20448 14924 20460
rect 14700 20420 14924 20448
rect 14700 20408 14706 20420
rect 14918 20408 14924 20420
rect 14976 20408 14982 20460
rect 15013 20451 15071 20457
rect 15013 20417 15025 20451
rect 15059 20448 15071 20451
rect 15102 20448 15108 20460
rect 15059 20420 15108 20448
rect 15059 20417 15071 20420
rect 15013 20411 15071 20417
rect 3513 20383 3571 20389
rect 3513 20349 3525 20383
rect 3559 20349 3571 20383
rect 3513 20343 3571 20349
rect 14277 20383 14335 20389
rect 14277 20349 14289 20383
rect 14323 20380 14335 20383
rect 15028 20380 15056 20411
rect 15102 20408 15108 20420
rect 15160 20408 15166 20460
rect 15197 20451 15255 20457
rect 15197 20417 15209 20451
rect 15243 20417 15255 20451
rect 15197 20411 15255 20417
rect 15289 20451 15347 20457
rect 15289 20417 15301 20451
rect 15335 20448 15347 20451
rect 15562 20448 15568 20460
rect 15335 20420 15568 20448
rect 15335 20417 15347 20420
rect 15289 20411 15347 20417
rect 14323 20352 15056 20380
rect 14323 20349 14335 20352
rect 14277 20343 14335 20349
rect 2866 20244 2872 20256
rect 2827 20216 2872 20244
rect 2866 20204 2872 20216
rect 2924 20204 2930 20256
rect 3528 20244 3556 20343
rect 13449 20315 13507 20321
rect 7576 20284 8524 20312
rect 3786 20244 3792 20256
rect 3528 20216 3792 20244
rect 3786 20204 3792 20216
rect 3844 20204 3850 20256
rect 4893 20247 4951 20253
rect 4893 20213 4905 20247
rect 4939 20244 4951 20247
rect 5537 20247 5595 20253
rect 5537 20244 5549 20247
rect 4939 20216 5549 20244
rect 4939 20213 4951 20216
rect 4893 20207 4951 20213
rect 5537 20213 5549 20216
rect 5583 20213 5595 20247
rect 6546 20244 6552 20256
rect 6507 20216 6552 20244
rect 5537 20207 5595 20213
rect 6546 20204 6552 20216
rect 6604 20204 6610 20256
rect 7576 20253 7604 20284
rect 7561 20247 7619 20253
rect 7561 20213 7573 20247
rect 7607 20213 7619 20247
rect 7561 20207 7619 20213
rect 7745 20247 7803 20253
rect 7745 20213 7757 20247
rect 7791 20244 7803 20247
rect 8386 20244 8392 20256
rect 7791 20216 8392 20244
rect 7791 20213 7803 20216
rect 7745 20207 7803 20213
rect 8386 20204 8392 20216
rect 8444 20204 8450 20256
rect 8496 20244 8524 20284
rect 13449 20281 13461 20315
rect 13495 20312 13507 20315
rect 15212 20312 15240 20411
rect 15562 20408 15568 20420
rect 15620 20408 15626 20460
rect 15856 20457 15884 20488
rect 16850 20476 16856 20488
rect 16908 20476 16914 20528
rect 16960 20516 16988 20556
rect 17681 20553 17693 20587
rect 17727 20584 17739 20587
rect 17770 20584 17776 20596
rect 17727 20556 17776 20584
rect 17727 20553 17739 20556
rect 17681 20547 17739 20553
rect 17770 20544 17776 20556
rect 17828 20544 17834 20596
rect 19797 20587 19855 20593
rect 19797 20553 19809 20587
rect 19843 20584 19855 20587
rect 20070 20584 20076 20596
rect 19843 20556 20076 20584
rect 19843 20553 19855 20556
rect 19797 20547 19855 20553
rect 20070 20544 20076 20556
rect 20128 20544 20134 20596
rect 24581 20587 24639 20593
rect 24581 20553 24593 20587
rect 24627 20584 24639 20587
rect 25406 20584 25412 20596
rect 24627 20556 25412 20584
rect 24627 20553 24639 20556
rect 24581 20547 24639 20553
rect 25406 20544 25412 20556
rect 25464 20544 25470 20596
rect 26878 20584 26884 20596
rect 26298 20556 26884 20584
rect 16960 20488 18736 20516
rect 15841 20451 15899 20457
rect 15841 20417 15853 20451
rect 15887 20417 15899 20451
rect 15841 20411 15899 20417
rect 15933 20451 15991 20457
rect 15933 20417 15945 20451
rect 15979 20448 15991 20451
rect 16482 20448 16488 20460
rect 15979 20420 16488 20448
rect 15979 20417 15991 20420
rect 15933 20411 15991 20417
rect 16482 20408 16488 20420
rect 16540 20408 16546 20460
rect 16669 20451 16727 20457
rect 16669 20417 16681 20451
rect 16715 20448 16727 20451
rect 16758 20448 16764 20460
rect 16715 20420 16764 20448
rect 16715 20417 16727 20420
rect 16669 20411 16727 20417
rect 16758 20408 16764 20420
rect 16816 20448 16822 20460
rect 16960 20448 16988 20488
rect 16816 20420 16988 20448
rect 17865 20451 17923 20457
rect 16816 20408 16822 20420
rect 17865 20417 17877 20451
rect 17911 20417 17923 20451
rect 17865 20411 17923 20417
rect 17880 20380 17908 20411
rect 17954 20408 17960 20460
rect 18012 20448 18018 20460
rect 18138 20448 18144 20460
rect 18012 20420 18057 20448
rect 18099 20420 18144 20448
rect 18012 20408 18018 20420
rect 18138 20408 18144 20420
rect 18196 20408 18202 20460
rect 18230 20408 18236 20460
rect 18288 20448 18294 20460
rect 18708 20457 18736 20488
rect 18782 20476 18788 20528
rect 18840 20516 18846 20528
rect 18877 20519 18935 20525
rect 18877 20516 18889 20519
rect 18840 20488 18889 20516
rect 18840 20476 18846 20488
rect 18877 20485 18889 20488
rect 18923 20485 18935 20519
rect 18877 20479 18935 20485
rect 18984 20488 20852 20516
rect 18693 20451 18751 20457
rect 18288 20420 18333 20448
rect 18288 20408 18294 20420
rect 18693 20417 18705 20451
rect 18739 20448 18751 20451
rect 18984 20448 19012 20488
rect 20070 20448 20076 20460
rect 18739 20420 19012 20448
rect 20031 20420 20076 20448
rect 18739 20417 18751 20420
rect 18693 20411 18751 20417
rect 20070 20408 20076 20420
rect 20128 20408 20134 20460
rect 20165 20451 20223 20457
rect 20165 20417 20177 20451
rect 20211 20417 20223 20451
rect 20165 20411 20223 20417
rect 18322 20380 18328 20392
rect 17880 20352 18328 20380
rect 18322 20340 18328 20352
rect 18380 20380 18386 20392
rect 18380 20352 19196 20380
rect 18380 20340 18386 20352
rect 16666 20312 16672 20324
rect 13495 20284 15148 20312
rect 15212 20284 16672 20312
rect 13495 20281 13507 20284
rect 13449 20275 13507 20281
rect 9953 20247 10011 20253
rect 9953 20244 9965 20247
rect 8496 20216 9965 20244
rect 9953 20213 9965 20216
rect 9999 20213 10011 20247
rect 15120 20244 15148 20284
rect 16666 20272 16672 20284
rect 16724 20272 16730 20324
rect 16022 20244 16028 20256
rect 15120 20216 16028 20244
rect 9953 20207 10011 20213
rect 16022 20204 16028 20216
rect 16080 20204 16086 20256
rect 16117 20247 16175 20253
rect 16117 20213 16129 20247
rect 16163 20244 16175 20247
rect 16574 20244 16580 20256
rect 16163 20216 16580 20244
rect 16163 20213 16175 20216
rect 16117 20207 16175 20213
rect 16574 20204 16580 20216
rect 16632 20204 16638 20256
rect 17034 20244 17040 20256
rect 16995 20216 17040 20244
rect 17034 20204 17040 20216
rect 17092 20204 17098 20256
rect 18414 20204 18420 20256
rect 18472 20244 18478 20256
rect 19061 20247 19119 20253
rect 19061 20244 19073 20247
rect 18472 20216 19073 20244
rect 18472 20204 18478 20216
rect 19061 20213 19073 20216
rect 19107 20213 19119 20247
rect 19168 20244 19196 20352
rect 20070 20272 20076 20324
rect 20128 20312 20134 20324
rect 20171 20312 20199 20411
rect 20254 20408 20260 20460
rect 20312 20448 20318 20460
rect 20438 20448 20444 20460
rect 20312 20420 20357 20448
rect 20399 20420 20444 20448
rect 20312 20408 20318 20420
rect 20438 20408 20444 20420
rect 20496 20408 20502 20460
rect 20824 20448 20852 20488
rect 20898 20476 20904 20528
rect 20956 20516 20962 20528
rect 20956 20488 22692 20516
rect 20956 20476 20962 20488
rect 22002 20448 22008 20460
rect 20824 20420 22008 20448
rect 22002 20408 22008 20420
rect 22060 20408 22066 20460
rect 22664 20457 22692 20488
rect 23566 20476 23572 20528
rect 23624 20516 23630 20528
rect 25501 20519 25559 20525
rect 25501 20516 25513 20519
rect 23624 20488 25513 20516
rect 23624 20476 23630 20488
rect 25501 20485 25513 20488
rect 25547 20485 25559 20519
rect 25501 20479 25559 20485
rect 22649 20451 22707 20457
rect 22649 20417 22661 20451
rect 22695 20417 22707 20451
rect 22649 20411 22707 20417
rect 22833 20451 22891 20457
rect 22833 20417 22845 20451
rect 22879 20448 22891 20451
rect 24486 20448 24492 20460
rect 22879 20420 24492 20448
rect 22879 20417 22891 20420
rect 22833 20411 22891 20417
rect 22664 20380 22692 20411
rect 24486 20408 24492 20420
rect 24544 20408 24550 20460
rect 24673 20451 24731 20457
rect 24673 20417 24685 20451
rect 24719 20417 24731 20451
rect 25130 20448 25136 20460
rect 25091 20420 25136 20448
rect 24673 20411 24731 20417
rect 24118 20380 24124 20392
rect 22664 20352 24124 20380
rect 24118 20340 24124 20352
rect 24176 20340 24182 20392
rect 24302 20340 24308 20392
rect 24360 20380 24366 20392
rect 24688 20380 24716 20411
rect 25130 20408 25136 20420
rect 25188 20408 25194 20460
rect 25222 20408 25228 20460
rect 25280 20448 25286 20460
rect 25406 20448 25412 20460
rect 25280 20420 25325 20448
rect 25367 20420 25412 20448
rect 25280 20408 25286 20420
rect 25406 20408 25412 20420
rect 25464 20408 25470 20460
rect 25639 20451 25697 20457
rect 25639 20417 25651 20451
rect 25685 20448 25697 20451
rect 26298 20448 26326 20556
rect 26878 20544 26884 20556
rect 26936 20584 26942 20596
rect 26936 20556 27384 20584
rect 26936 20544 26942 20556
rect 26973 20519 27031 20525
rect 26973 20485 26985 20519
rect 27019 20516 27031 20519
rect 27246 20516 27252 20528
rect 27019 20488 27252 20516
rect 27019 20485 27031 20488
rect 26973 20479 27031 20485
rect 27246 20476 27252 20488
rect 27304 20476 27310 20528
rect 27356 20516 27384 20556
rect 27798 20544 27804 20596
rect 27856 20584 27862 20596
rect 27893 20587 27951 20593
rect 27893 20584 27905 20587
rect 27856 20556 27905 20584
rect 27856 20544 27862 20556
rect 27893 20553 27905 20556
rect 27939 20553 27951 20587
rect 27893 20547 27951 20553
rect 28445 20587 28503 20593
rect 28445 20553 28457 20587
rect 28491 20584 28503 20587
rect 28718 20584 28724 20596
rect 28491 20556 28724 20584
rect 28491 20553 28503 20556
rect 28445 20547 28503 20553
rect 28718 20544 28724 20556
rect 28776 20544 28782 20596
rect 28810 20544 28816 20596
rect 28868 20544 28874 20596
rect 28994 20544 29000 20596
rect 29052 20584 29058 20596
rect 29914 20584 29920 20596
rect 29052 20556 29920 20584
rect 29052 20544 29058 20556
rect 29914 20544 29920 20556
rect 29972 20584 29978 20596
rect 30190 20584 30196 20596
rect 29972 20556 30196 20584
rect 29972 20544 29978 20556
rect 30190 20544 30196 20556
rect 30248 20544 30254 20596
rect 28350 20516 28356 20528
rect 27356 20488 28356 20516
rect 28350 20476 28356 20488
rect 28408 20476 28414 20528
rect 25685 20420 26326 20448
rect 27157 20451 27215 20457
rect 25685 20417 25697 20420
rect 25639 20411 25697 20417
rect 27157 20417 27169 20451
rect 27203 20448 27215 20451
rect 27798 20448 27804 20460
rect 27203 20420 27804 20448
rect 27203 20417 27215 20420
rect 27157 20411 27215 20417
rect 24360 20352 24716 20380
rect 24360 20340 24366 20352
rect 24854 20340 24860 20392
rect 24912 20380 24918 20392
rect 25654 20380 25682 20411
rect 27798 20408 27804 20420
rect 27856 20408 27862 20460
rect 27985 20451 28043 20457
rect 27985 20417 27997 20451
rect 28031 20448 28043 20451
rect 28074 20448 28080 20460
rect 28031 20420 28080 20448
rect 28031 20417 28043 20420
rect 27985 20411 28043 20417
rect 28074 20408 28080 20420
rect 28132 20408 28138 20460
rect 28828 20457 28856 20544
rect 29822 20525 29828 20528
rect 29816 20516 29828 20525
rect 29783 20488 29828 20516
rect 29816 20479 29828 20488
rect 29822 20476 29828 20479
rect 29880 20476 29886 20528
rect 28721 20451 28779 20457
rect 28700 20417 28733 20451
rect 28767 20417 28779 20451
rect 28700 20411 28779 20417
rect 28813 20451 28871 20457
rect 28813 20417 28825 20451
rect 28859 20417 28871 20451
rect 28813 20411 28871 20417
rect 24912 20352 25682 20380
rect 24912 20340 24918 20352
rect 26694 20340 26700 20392
rect 26752 20380 26758 20392
rect 28700 20380 28728 20411
rect 28902 20408 28908 20460
rect 28960 20448 28966 20460
rect 29089 20451 29147 20457
rect 28960 20420 29005 20448
rect 28960 20408 28966 20420
rect 29089 20417 29101 20451
rect 29135 20448 29147 20451
rect 30742 20448 30748 20460
rect 29135 20420 30748 20448
rect 29135 20417 29147 20420
rect 29089 20411 29147 20417
rect 30742 20408 30748 20420
rect 30800 20408 30806 20460
rect 31754 20408 31760 20460
rect 31812 20448 31818 20460
rect 32493 20451 32551 20457
rect 32493 20448 32505 20451
rect 31812 20420 32505 20448
rect 31812 20408 31818 20420
rect 32493 20417 32505 20420
rect 32539 20417 32551 20451
rect 32493 20411 32551 20417
rect 33870 20408 33876 20460
rect 33928 20448 33934 20460
rect 33965 20451 34023 20457
rect 33965 20448 33977 20451
rect 33928 20420 33977 20448
rect 33928 20408 33934 20420
rect 33965 20417 33977 20420
rect 34011 20417 34023 20451
rect 33965 20411 34023 20417
rect 34514 20408 34520 20460
rect 34572 20448 34578 20460
rect 34885 20451 34943 20457
rect 34885 20448 34897 20451
rect 34572 20420 34897 20448
rect 34572 20408 34578 20420
rect 34885 20417 34897 20420
rect 34931 20417 34943 20451
rect 34885 20411 34943 20417
rect 29362 20380 29368 20392
rect 26752 20352 29368 20380
rect 26752 20340 26758 20352
rect 29362 20340 29368 20352
rect 29420 20340 29426 20392
rect 29549 20383 29607 20389
rect 29549 20349 29561 20383
rect 29595 20349 29607 20383
rect 29549 20343 29607 20349
rect 32769 20383 32827 20389
rect 32769 20349 32781 20383
rect 32815 20380 32827 20383
rect 33686 20380 33692 20392
rect 32815 20352 33692 20380
rect 32815 20349 32827 20352
rect 32769 20343 32827 20349
rect 20128 20284 20199 20312
rect 20128 20272 20134 20284
rect 21726 20272 21732 20324
rect 21784 20312 21790 20324
rect 21784 20284 28580 20312
rect 21784 20272 21790 20284
rect 21082 20244 21088 20256
rect 19168 20216 21088 20244
rect 19061 20207 19119 20213
rect 21082 20204 21088 20216
rect 21140 20204 21146 20256
rect 23017 20247 23075 20253
rect 23017 20213 23029 20247
rect 23063 20244 23075 20247
rect 23474 20244 23480 20256
rect 23063 20216 23480 20244
rect 23063 20213 23075 20216
rect 23017 20207 23075 20213
rect 23474 20204 23480 20216
rect 23532 20204 23538 20256
rect 23750 20204 23756 20256
rect 23808 20244 23814 20256
rect 24670 20244 24676 20256
rect 23808 20216 24676 20244
rect 23808 20204 23814 20216
rect 24670 20204 24676 20216
rect 24728 20204 24734 20256
rect 25777 20247 25835 20253
rect 25777 20213 25789 20247
rect 25823 20244 25835 20247
rect 26510 20244 26516 20256
rect 25823 20216 26516 20244
rect 25823 20213 25835 20216
rect 25777 20207 25835 20213
rect 26510 20204 26516 20216
rect 26568 20204 26574 20256
rect 26970 20204 26976 20256
rect 27028 20244 27034 20256
rect 27341 20247 27399 20253
rect 27341 20244 27353 20247
rect 27028 20216 27353 20244
rect 27028 20204 27034 20216
rect 27341 20213 27353 20216
rect 27387 20213 27399 20247
rect 28552 20244 28580 20284
rect 28718 20272 28724 20324
rect 28776 20312 28782 20324
rect 29564 20312 29592 20343
rect 33686 20340 33692 20352
rect 33744 20340 33750 20392
rect 34241 20383 34299 20389
rect 34241 20349 34253 20383
rect 34287 20380 34299 20383
rect 34790 20380 34796 20392
rect 34287 20352 34796 20380
rect 34287 20349 34299 20352
rect 34241 20343 34299 20349
rect 34790 20340 34796 20352
rect 34848 20340 34854 20392
rect 28776 20284 29592 20312
rect 28776 20272 28782 20284
rect 31294 20272 31300 20324
rect 31352 20312 31358 20324
rect 32677 20315 32735 20321
rect 32677 20312 32689 20315
rect 31352 20284 32689 20312
rect 31352 20272 31358 20284
rect 32677 20281 32689 20284
rect 32723 20312 32735 20315
rect 32858 20312 32864 20324
rect 32723 20284 32864 20312
rect 32723 20281 32735 20284
rect 32677 20275 32735 20281
rect 32858 20272 32864 20284
rect 32916 20312 32922 20324
rect 34149 20315 34207 20321
rect 34149 20312 34161 20315
rect 32916 20284 34161 20312
rect 32916 20272 32922 20284
rect 34149 20281 34161 20284
rect 34195 20281 34207 20315
rect 34149 20275 34207 20281
rect 28994 20244 29000 20256
rect 28552 20216 29000 20244
rect 27341 20207 27399 20213
rect 28994 20204 29000 20216
rect 29052 20204 29058 20256
rect 29362 20204 29368 20256
rect 29420 20244 29426 20256
rect 30926 20244 30932 20256
rect 29420 20216 30932 20244
rect 29420 20204 29426 20216
rect 30926 20204 30932 20216
rect 30984 20204 30990 20256
rect 32306 20244 32312 20256
rect 32267 20216 32312 20244
rect 32306 20204 32312 20216
rect 32364 20204 32370 20256
rect 33134 20204 33140 20256
rect 33192 20244 33198 20256
rect 33781 20247 33839 20253
rect 33781 20244 33793 20247
rect 33192 20216 33793 20244
rect 33192 20204 33198 20216
rect 33781 20213 33793 20216
rect 33827 20213 33839 20247
rect 33781 20207 33839 20213
rect 34330 20204 34336 20256
rect 34388 20244 34394 20256
rect 34701 20247 34759 20253
rect 34701 20244 34713 20247
rect 34388 20216 34713 20244
rect 34388 20204 34394 20216
rect 34701 20213 34713 20216
rect 34747 20213 34759 20247
rect 34701 20207 34759 20213
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 5169 20043 5227 20049
rect 5169 20009 5181 20043
rect 5215 20040 5227 20043
rect 6546 20040 6552 20052
rect 5215 20012 6552 20040
rect 5215 20009 5227 20012
rect 5169 20003 5227 20009
rect 6546 20000 6552 20012
rect 6604 20000 6610 20052
rect 7561 20043 7619 20049
rect 7561 20009 7573 20043
rect 7607 20009 7619 20043
rect 7561 20003 7619 20009
rect 8205 20043 8263 20049
rect 8205 20009 8217 20043
rect 8251 20040 8263 20043
rect 8662 20040 8668 20052
rect 8251 20012 8668 20040
rect 8251 20009 8263 20012
rect 8205 20003 8263 20009
rect 2866 19864 2872 19916
rect 2924 19904 2930 19916
rect 7576 19904 7604 20003
rect 8662 20000 8668 20012
rect 8720 20000 8726 20052
rect 10321 20043 10379 20049
rect 10321 20040 10333 20043
rect 8772 20012 10333 20040
rect 7745 19975 7803 19981
rect 7745 19941 7757 19975
rect 7791 19972 7803 19975
rect 8478 19972 8484 19984
rect 7791 19944 8484 19972
rect 7791 19941 7803 19944
rect 7745 19935 7803 19941
rect 8478 19932 8484 19944
rect 8536 19932 8542 19984
rect 8772 19904 8800 20012
rect 10321 20009 10333 20012
rect 10367 20009 10379 20043
rect 10321 20003 10379 20009
rect 17310 20000 17316 20052
rect 17368 20040 17374 20052
rect 17368 20012 19932 20040
rect 17368 20000 17374 20012
rect 14550 19932 14556 19984
rect 14608 19972 14614 19984
rect 15562 19972 15568 19984
rect 14608 19944 15568 19972
rect 14608 19932 14614 19944
rect 15562 19932 15568 19944
rect 15620 19932 15626 19984
rect 18322 19932 18328 19984
rect 18380 19932 18386 19984
rect 8938 19904 8944 19916
rect 2924 19876 3924 19904
rect 7576 19876 8800 19904
rect 8899 19876 8944 19904
rect 2924 19864 2930 19876
rect 3786 19836 3792 19848
rect 3747 19808 3792 19836
rect 3786 19796 3792 19808
rect 3844 19796 3850 19848
rect 3896 19836 3924 19876
rect 8938 19864 8944 19876
rect 8996 19864 9002 19916
rect 4045 19839 4103 19845
rect 4045 19836 4057 19839
rect 3896 19808 4057 19836
rect 4045 19805 4057 19808
rect 4091 19805 4103 19839
rect 6914 19836 6920 19848
rect 6875 19808 6920 19836
rect 4045 19799 4103 19805
rect 6914 19796 6920 19808
rect 6972 19796 6978 19848
rect 8386 19836 8392 19848
rect 8347 19808 8392 19836
rect 8386 19796 8392 19808
rect 8444 19796 8450 19848
rect 9030 19796 9036 19848
rect 9088 19836 9094 19848
rect 9197 19839 9255 19845
rect 9197 19836 9209 19839
rect 9088 19808 9209 19836
rect 9088 19796 9094 19808
rect 9197 19805 9209 19808
rect 9243 19805 9255 19839
rect 9197 19799 9255 19805
rect 10870 19796 10876 19848
rect 10928 19836 10934 19848
rect 10965 19839 11023 19845
rect 10965 19836 10977 19839
rect 10928 19808 10977 19836
rect 10928 19796 10934 19808
rect 10965 19805 10977 19808
rect 11011 19805 11023 19839
rect 10965 19799 11023 19805
rect 15194 19796 15200 19848
rect 15252 19836 15258 19848
rect 15580 19845 15608 19932
rect 15473 19839 15531 19845
rect 15473 19836 15485 19839
rect 15252 19808 15485 19836
rect 15252 19796 15258 19808
rect 15473 19805 15485 19808
rect 15519 19805 15531 19839
rect 15473 19799 15531 19805
rect 15565 19839 15623 19845
rect 15565 19805 15577 19839
rect 15611 19805 15623 19839
rect 15565 19799 15623 19805
rect 15657 19839 15715 19845
rect 15657 19805 15669 19839
rect 15703 19805 15715 19839
rect 15657 19799 15715 19805
rect 15841 19839 15899 19845
rect 15841 19805 15853 19839
rect 15887 19805 15899 19839
rect 15841 19799 15899 19805
rect 7374 19768 7380 19780
rect 7287 19740 7380 19768
rect 7374 19728 7380 19740
rect 7432 19728 7438 19780
rect 7558 19728 7564 19780
rect 7616 19777 7622 19780
rect 7616 19771 7635 19777
rect 7623 19737 7635 19771
rect 7616 19731 7635 19737
rect 7616 19728 7622 19731
rect 11054 19728 11060 19780
rect 11112 19768 11118 19780
rect 11210 19771 11268 19777
rect 11210 19768 11222 19771
rect 11112 19740 11222 19768
rect 11112 19728 11118 19740
rect 11210 19737 11222 19740
rect 11256 19737 11268 19771
rect 11210 19731 11268 19737
rect 11698 19728 11704 19780
rect 11756 19768 11762 19780
rect 13998 19768 14004 19780
rect 11756 19740 14004 19768
rect 11756 19728 11762 19740
rect 13998 19728 14004 19740
rect 14056 19768 14062 19780
rect 14093 19771 14151 19777
rect 14093 19768 14105 19771
rect 14056 19740 14105 19768
rect 14056 19728 14062 19740
rect 14093 19737 14105 19740
rect 14139 19737 14151 19771
rect 14274 19768 14280 19780
rect 14235 19740 14280 19768
rect 14093 19731 14151 19737
rect 14274 19728 14280 19740
rect 14332 19728 14338 19780
rect 15672 19768 15700 19799
rect 14476 19740 15700 19768
rect 15856 19768 15884 19799
rect 16298 19796 16304 19848
rect 16356 19836 16362 19848
rect 16853 19839 16911 19845
rect 16853 19836 16865 19839
rect 16356 19808 16865 19836
rect 16356 19796 16362 19808
rect 16853 19805 16865 19808
rect 16899 19805 16911 19839
rect 18230 19836 18236 19848
rect 18191 19808 18236 19836
rect 16853 19799 16911 19805
rect 18230 19796 18236 19808
rect 18288 19796 18294 19848
rect 18340 19845 18368 19932
rect 19904 19913 19932 20012
rect 20622 20000 20628 20052
rect 20680 20040 20686 20052
rect 20806 20040 20812 20052
rect 20680 20012 20812 20040
rect 20680 20000 20686 20012
rect 20806 20000 20812 20012
rect 20864 20000 20870 20052
rect 23382 20000 23388 20052
rect 23440 20040 23446 20052
rect 25222 20040 25228 20052
rect 23440 20012 25228 20040
rect 23440 20000 23446 20012
rect 19889 19907 19947 19913
rect 19889 19873 19901 19907
rect 19935 19873 19947 19907
rect 21726 19904 21732 19916
rect 21687 19876 21732 19904
rect 19889 19867 19947 19873
rect 18322 19839 18380 19845
rect 18322 19805 18334 19839
rect 18368 19805 18380 19839
rect 18322 19799 18380 19805
rect 18414 19796 18420 19848
rect 18472 19836 18478 19848
rect 18601 19839 18659 19845
rect 18472 19808 18517 19836
rect 18472 19796 18478 19808
rect 18601 19805 18613 19839
rect 18647 19836 18659 19839
rect 18690 19836 18696 19848
rect 18647 19808 18696 19836
rect 18647 19805 18659 19808
rect 18601 19799 18659 19805
rect 18690 19796 18696 19808
rect 18748 19796 18754 19848
rect 19904 19836 19932 19867
rect 21726 19864 21732 19876
rect 21784 19864 21790 19916
rect 22002 19864 22008 19916
rect 22060 19904 22066 19916
rect 22060 19876 22105 19904
rect 22060 19864 22066 19876
rect 23198 19864 23204 19916
rect 23256 19904 23262 19916
rect 23566 19904 23572 19916
rect 23256 19876 23572 19904
rect 23256 19864 23262 19876
rect 20438 19836 20444 19848
rect 19904 19808 20444 19836
rect 20438 19796 20444 19808
rect 20496 19796 20502 19848
rect 22646 19796 22652 19848
rect 22704 19836 22710 19848
rect 23400 19845 23428 19876
rect 23566 19864 23572 19876
rect 23624 19864 23630 19916
rect 23293 19839 23351 19845
rect 23293 19836 23305 19839
rect 22704 19808 23305 19836
rect 22704 19796 22710 19808
rect 23293 19805 23305 19808
rect 23339 19805 23351 19839
rect 23293 19799 23351 19805
rect 23385 19839 23443 19845
rect 23385 19805 23397 19839
rect 23431 19805 23443 19839
rect 23385 19799 23443 19805
rect 23474 19796 23480 19848
rect 23532 19836 23538 19848
rect 23676 19845 23704 20012
rect 25222 20000 25228 20012
rect 25280 20000 25286 20052
rect 30558 20000 30564 20052
rect 30616 20040 30622 20052
rect 31389 20043 31447 20049
rect 31389 20040 31401 20043
rect 30616 20012 31401 20040
rect 30616 20000 30622 20012
rect 31389 20009 31401 20012
rect 31435 20009 31447 20043
rect 33686 20040 33692 20052
rect 33647 20012 33692 20040
rect 31389 20003 31447 20009
rect 25130 19972 25136 19984
rect 24412 19944 25136 19972
rect 24412 19845 24440 19944
rect 25130 19932 25136 19944
rect 25188 19932 25194 19984
rect 27706 19972 27712 19984
rect 27632 19944 27712 19972
rect 24670 19864 24676 19916
rect 24728 19864 24734 19916
rect 23661 19839 23719 19845
rect 23532 19808 23577 19836
rect 23532 19796 23538 19808
rect 23661 19805 23673 19839
rect 23707 19805 23719 19839
rect 23661 19799 23719 19805
rect 24397 19839 24455 19845
rect 24397 19805 24409 19839
rect 24443 19805 24455 19839
rect 24397 19799 24455 19805
rect 24486 19796 24492 19848
rect 24544 19836 24550 19848
rect 24688 19836 24716 19864
rect 24544 19808 24589 19836
rect 24688 19808 24808 19836
rect 24544 19796 24550 19808
rect 16390 19768 16396 19780
rect 15856 19740 16396 19768
rect 6454 19660 6460 19712
rect 6512 19700 6518 19712
rect 6733 19703 6791 19709
rect 6733 19700 6745 19703
rect 6512 19672 6745 19700
rect 6512 19660 6518 19672
rect 6733 19669 6745 19672
rect 6779 19700 6791 19703
rect 7392 19700 7420 19728
rect 12342 19700 12348 19712
rect 6779 19672 7420 19700
rect 12303 19672 12348 19700
rect 6779 19669 6791 19672
rect 6733 19663 6791 19669
rect 12342 19660 12348 19672
rect 12400 19660 12406 19712
rect 13814 19660 13820 19712
rect 13872 19700 13878 19712
rect 14476 19709 14504 19740
rect 16390 19728 16396 19740
rect 16448 19728 16454 19780
rect 16669 19771 16727 19777
rect 16669 19737 16681 19771
rect 16715 19768 16727 19771
rect 16758 19768 16764 19780
rect 16715 19740 16764 19768
rect 16715 19737 16727 19740
rect 16669 19731 16727 19737
rect 16758 19728 16764 19740
rect 16816 19728 16822 19780
rect 20162 19777 20168 19780
rect 20156 19731 20168 19777
rect 20220 19768 20226 19780
rect 20220 19740 20256 19768
rect 20162 19728 20168 19731
rect 20220 19728 20226 19740
rect 23750 19728 23756 19780
rect 23808 19768 23814 19780
rect 24504 19768 24532 19796
rect 24780 19777 24808 19808
rect 24854 19796 24860 19848
rect 24912 19845 24918 19848
rect 24912 19836 24920 19845
rect 24912 19808 24957 19836
rect 24912 19799 24920 19808
rect 24912 19796 24918 19799
rect 25130 19796 25136 19848
rect 25188 19836 25194 19848
rect 26329 19839 26387 19845
rect 26329 19836 26341 19839
rect 25188 19808 26341 19836
rect 25188 19796 25194 19808
rect 26329 19805 26341 19808
rect 26375 19805 26387 19839
rect 26329 19799 26387 19805
rect 26477 19839 26535 19845
rect 26477 19805 26489 19839
rect 26523 19836 26535 19839
rect 26694 19836 26700 19848
rect 26523 19805 26556 19836
rect 26655 19808 26700 19836
rect 26477 19799 26556 19805
rect 23808 19740 24532 19768
rect 24673 19771 24731 19777
rect 23808 19728 23814 19740
rect 24673 19737 24685 19771
rect 24719 19737 24731 19771
rect 24673 19731 24731 19737
rect 24765 19771 24823 19777
rect 24765 19737 24777 19771
rect 24811 19737 24823 19771
rect 25406 19768 25412 19780
rect 24765 19731 24823 19737
rect 24872 19740 25412 19768
rect 14461 19703 14519 19709
rect 14461 19700 14473 19703
rect 13872 19672 14473 19700
rect 13872 19660 13878 19672
rect 14461 19669 14473 19672
rect 14507 19669 14519 19703
rect 15194 19700 15200 19712
rect 15155 19672 15200 19700
rect 14461 19663 14519 19669
rect 15194 19660 15200 19672
rect 15252 19660 15258 19712
rect 16574 19660 16580 19712
rect 16632 19700 16638 19712
rect 17037 19703 17095 19709
rect 17037 19700 17049 19703
rect 16632 19672 17049 19700
rect 16632 19660 16638 19672
rect 17037 19669 17049 19672
rect 17083 19669 17095 19703
rect 17037 19663 17095 19669
rect 17957 19703 18015 19709
rect 17957 19669 17969 19703
rect 18003 19700 18015 19703
rect 18414 19700 18420 19712
rect 18003 19672 18420 19700
rect 18003 19669 18015 19672
rect 17957 19663 18015 19669
rect 18414 19660 18420 19672
rect 18472 19660 18478 19712
rect 21269 19703 21327 19709
rect 21269 19669 21281 19703
rect 21315 19700 21327 19703
rect 22370 19700 22376 19712
rect 21315 19672 22376 19700
rect 21315 19669 21327 19672
rect 21269 19663 21327 19669
rect 22370 19660 22376 19672
rect 22428 19660 22434 19712
rect 23014 19700 23020 19712
rect 22975 19672 23020 19700
rect 23014 19660 23020 19672
rect 23072 19660 23078 19712
rect 24688 19700 24716 19731
rect 24872 19700 24900 19740
rect 25406 19728 25412 19740
rect 25464 19728 25470 19780
rect 24688 19672 24900 19700
rect 24946 19660 24952 19712
rect 25004 19700 25010 19712
rect 25041 19703 25099 19709
rect 25041 19700 25053 19703
rect 25004 19672 25053 19700
rect 25004 19660 25010 19672
rect 25041 19669 25053 19672
rect 25087 19669 25099 19703
rect 26528 19700 26556 19799
rect 26694 19796 26700 19808
rect 26752 19796 26758 19848
rect 26878 19845 26884 19848
rect 26835 19839 26884 19845
rect 26835 19805 26847 19839
rect 26881 19805 26884 19839
rect 26835 19799 26884 19805
rect 26878 19796 26884 19799
rect 26936 19796 26942 19848
rect 27430 19836 27436 19848
rect 26988 19808 27436 19836
rect 26605 19771 26663 19777
rect 26605 19737 26617 19771
rect 26651 19768 26663 19771
rect 26988 19768 27016 19808
rect 27430 19796 27436 19808
rect 27488 19796 27494 19848
rect 27632 19833 27660 19944
rect 27706 19932 27712 19944
rect 27764 19972 27770 19984
rect 28166 19972 28172 19984
rect 27764 19944 28172 19972
rect 27764 19932 27770 19944
rect 28166 19932 28172 19944
rect 28224 19932 28230 19984
rect 28994 19932 29000 19984
rect 29052 19972 29058 19984
rect 31294 19972 31300 19984
rect 29052 19944 31300 19972
rect 29052 19932 29058 19944
rect 31294 19932 31300 19944
rect 31352 19932 31358 19984
rect 28442 19864 28448 19916
rect 28500 19904 28506 19916
rect 31404 19904 31432 20003
rect 33686 20000 33692 20012
rect 33744 20000 33750 20052
rect 32309 19907 32367 19913
rect 32309 19904 32321 19907
rect 28500 19876 30144 19904
rect 31404 19876 32321 19904
rect 28500 19864 28506 19876
rect 27689 19839 27747 19845
rect 27689 19833 27701 19839
rect 27632 19805 27701 19833
rect 27735 19805 27747 19839
rect 27801 19839 27859 19845
rect 27801 19833 27813 19839
rect 27689 19799 27747 19805
rect 27797 19805 27813 19833
rect 27847 19805 27859 19839
rect 27797 19799 27859 19805
rect 26651 19740 27016 19768
rect 27797 19768 27825 19799
rect 27890 19796 27896 19848
rect 27948 19836 27954 19848
rect 28077 19839 28135 19845
rect 27948 19808 27993 19836
rect 27948 19796 27954 19808
rect 28077 19805 28089 19839
rect 28123 19836 28135 19839
rect 28166 19836 28172 19848
rect 28123 19808 28172 19836
rect 28123 19805 28135 19808
rect 28077 19799 28135 19805
rect 28166 19796 28172 19808
rect 28224 19796 28230 19848
rect 30116 19845 30144 19876
rect 32309 19873 32321 19876
rect 32355 19873 32367 19907
rect 32309 19867 32367 19873
rect 33778 19864 33784 19916
rect 33836 19904 33842 19916
rect 33836 19876 34928 19904
rect 33836 19864 33842 19876
rect 30101 19839 30159 19845
rect 30101 19805 30113 19839
rect 30147 19805 30159 19839
rect 30101 19799 30159 19805
rect 32950 19796 32956 19848
rect 33008 19836 33014 19848
rect 34900 19845 34928 19876
rect 34701 19839 34759 19845
rect 34701 19836 34713 19839
rect 33008 19808 34713 19836
rect 33008 19796 33014 19808
rect 34701 19805 34713 19808
rect 34747 19805 34759 19839
rect 34701 19799 34759 19805
rect 34885 19839 34943 19845
rect 34885 19805 34897 19839
rect 34931 19805 34943 19839
rect 34885 19799 34943 19805
rect 28350 19768 28356 19780
rect 27797 19740 28356 19768
rect 26651 19737 26663 19740
rect 26605 19731 26663 19737
rect 28350 19728 28356 19740
rect 28408 19728 28414 19780
rect 32214 19728 32220 19780
rect 32272 19768 32278 19780
rect 32554 19771 32612 19777
rect 32554 19768 32566 19771
rect 32272 19740 32566 19768
rect 32272 19728 32278 19740
rect 32554 19737 32566 19740
rect 32600 19737 32612 19771
rect 32554 19731 32612 19737
rect 26694 19700 26700 19712
rect 26528 19672 26700 19700
rect 25041 19663 25099 19669
rect 26694 19660 26700 19672
rect 26752 19660 26758 19712
rect 26973 19703 27031 19709
rect 26973 19669 26985 19703
rect 27019 19700 27031 19703
rect 27154 19700 27160 19712
rect 27019 19672 27160 19700
rect 27019 19669 27031 19672
rect 26973 19663 27031 19669
rect 27154 19660 27160 19672
rect 27212 19660 27218 19712
rect 27430 19700 27436 19712
rect 27391 19672 27436 19700
rect 27430 19660 27436 19672
rect 27488 19660 27494 19712
rect 35069 19703 35127 19709
rect 35069 19669 35081 19703
rect 35115 19700 35127 19703
rect 37274 19700 37280 19712
rect 35115 19672 37280 19700
rect 35115 19669 35127 19672
rect 35069 19663 35127 19669
rect 37274 19660 37280 19672
rect 37332 19660 37338 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 4985 19499 5043 19505
rect 4985 19465 4997 19499
rect 5031 19496 5043 19499
rect 5074 19496 5080 19508
rect 5031 19468 5080 19496
rect 5031 19465 5043 19468
rect 4985 19459 5043 19465
rect 5074 19456 5080 19468
rect 5132 19456 5138 19508
rect 5629 19499 5687 19505
rect 5629 19465 5641 19499
rect 5675 19496 5687 19499
rect 5675 19468 6500 19496
rect 5675 19465 5687 19468
rect 5629 19459 5687 19465
rect 4617 19431 4675 19437
rect 4617 19397 4629 19431
rect 4663 19397 4675 19431
rect 4617 19391 4675 19397
rect 4833 19431 4891 19437
rect 4833 19397 4845 19431
rect 4879 19428 4891 19431
rect 5350 19428 5356 19440
rect 4879 19400 5356 19428
rect 4879 19397 4891 19400
rect 4833 19391 4891 19397
rect 4632 19360 4660 19391
rect 5350 19388 5356 19400
rect 5408 19388 5414 19440
rect 5534 19388 5540 19440
rect 5592 19428 5598 19440
rect 6472 19428 6500 19468
rect 9490 19456 9496 19508
rect 9548 19496 9554 19508
rect 9953 19499 10011 19505
rect 9953 19496 9965 19499
rect 9548 19468 9965 19496
rect 9548 19456 9554 19468
rect 9953 19465 9965 19468
rect 9999 19465 10011 19499
rect 9953 19459 10011 19465
rect 10870 19456 10876 19508
rect 10928 19496 10934 19508
rect 13173 19499 13231 19505
rect 13173 19496 13185 19499
rect 10928 19468 13185 19496
rect 10928 19456 10934 19468
rect 13173 19465 13185 19468
rect 13219 19465 13231 19499
rect 13173 19459 13231 19465
rect 6610 19431 6668 19437
rect 6610 19428 6622 19431
rect 5592 19400 6408 19428
rect 6472 19400 6622 19428
rect 5592 19388 5598 19400
rect 5626 19360 5632 19372
rect 4632 19332 5632 19360
rect 5626 19320 5632 19332
rect 5684 19320 5690 19372
rect 5810 19360 5816 19372
rect 5771 19332 5816 19360
rect 5810 19320 5816 19332
rect 5868 19320 5874 19372
rect 6380 19369 6408 19400
rect 6610 19397 6622 19400
rect 6656 19397 6668 19431
rect 8938 19428 8944 19440
rect 6610 19391 6668 19397
rect 8588 19400 8944 19428
rect 8588 19369 8616 19400
rect 8938 19388 8944 19400
rect 8996 19388 9002 19440
rect 9214 19388 9220 19440
rect 9272 19428 9278 19440
rect 11885 19431 11943 19437
rect 11885 19428 11897 19431
rect 9272 19400 11897 19428
rect 9272 19388 9278 19400
rect 11885 19397 11897 19400
rect 11931 19397 11943 19431
rect 11885 19391 11943 19397
rect 6365 19363 6423 19369
rect 6365 19329 6377 19363
rect 6411 19329 6423 19363
rect 6365 19323 6423 19329
rect 8573 19363 8631 19369
rect 8573 19329 8585 19363
rect 8619 19329 8631 19363
rect 8573 19323 8631 19329
rect 8662 19320 8668 19372
rect 8720 19360 8726 19372
rect 8829 19363 8887 19369
rect 8829 19360 8841 19363
rect 8720 19332 8841 19360
rect 8720 19320 8726 19332
rect 8829 19329 8841 19332
rect 8875 19329 8887 19363
rect 8829 19323 8887 19329
rect 10597 19363 10655 19369
rect 10597 19329 10609 19363
rect 10643 19329 10655 19363
rect 10778 19360 10784 19372
rect 10739 19332 10784 19360
rect 10597 19323 10655 19329
rect 10612 19292 10640 19323
rect 10778 19320 10784 19332
rect 10836 19320 10842 19372
rect 13188 19360 13216 19459
rect 14274 19456 14280 19508
rect 14332 19496 14338 19508
rect 15473 19499 15531 19505
rect 15473 19496 15485 19499
rect 14332 19468 15485 19496
rect 14332 19456 14338 19468
rect 15473 19465 15485 19468
rect 15519 19465 15531 19499
rect 15473 19459 15531 19465
rect 16758 19456 16764 19508
rect 16816 19496 16822 19508
rect 17126 19496 17132 19508
rect 16816 19468 17132 19496
rect 16816 19456 16822 19468
rect 17126 19456 17132 19468
rect 17184 19456 17190 19508
rect 18693 19499 18751 19505
rect 18693 19465 18705 19499
rect 18739 19496 18751 19499
rect 20438 19496 20444 19508
rect 18739 19468 19104 19496
rect 20399 19468 20444 19496
rect 18739 19465 18751 19468
rect 18693 19459 18751 19465
rect 14360 19431 14418 19437
rect 14360 19397 14372 19431
rect 14406 19428 14418 19431
rect 15194 19428 15200 19440
rect 14406 19400 15200 19428
rect 14406 19397 14418 19400
rect 14360 19391 14418 19397
rect 15194 19388 15200 19400
rect 15252 19388 15258 19440
rect 17954 19428 17960 19440
rect 16132 19400 16896 19428
rect 14093 19363 14151 19369
rect 14093 19360 14105 19363
rect 13188 19332 14105 19360
rect 14093 19329 14105 19332
rect 14139 19329 14151 19363
rect 15930 19360 15936 19372
rect 15891 19332 15936 19360
rect 14093 19323 14151 19329
rect 15930 19320 15936 19332
rect 15988 19320 15994 19372
rect 16022 19320 16028 19372
rect 16080 19360 16086 19372
rect 16132 19369 16160 19400
rect 16868 19369 16896 19400
rect 17144 19400 17960 19428
rect 16117 19363 16175 19369
rect 16117 19360 16129 19363
rect 16080 19332 16129 19360
rect 16080 19320 16086 19332
rect 16117 19329 16129 19332
rect 16163 19329 16175 19363
rect 16117 19323 16175 19329
rect 16669 19363 16727 19369
rect 16669 19329 16681 19363
rect 16715 19360 16727 19363
rect 16853 19363 16911 19369
rect 16715 19332 16804 19360
rect 16715 19329 16727 19332
rect 16669 19323 16727 19329
rect 11698 19292 11704 19304
rect 10612 19264 11704 19292
rect 11698 19252 11704 19264
rect 11756 19252 11762 19304
rect 16776 19292 16804 19332
rect 16853 19329 16865 19363
rect 16899 19329 16911 19363
rect 17144 19360 17172 19400
rect 17954 19388 17960 19400
rect 18012 19388 18018 19440
rect 18230 19388 18236 19440
rect 18288 19428 18294 19440
rect 18966 19428 18972 19440
rect 18288 19400 18972 19428
rect 18288 19388 18294 19400
rect 18966 19388 18972 19400
rect 19024 19388 19030 19440
rect 17310 19360 17316 19372
rect 16853 19323 16911 19329
rect 16960 19332 17172 19360
rect 17271 19332 17316 19360
rect 16960 19292 16988 19332
rect 17310 19320 17316 19332
rect 17368 19320 17374 19372
rect 17580 19363 17638 19369
rect 17580 19329 17592 19363
rect 17626 19360 17638 19363
rect 17862 19360 17868 19372
rect 17626 19332 17868 19360
rect 17626 19329 17638 19332
rect 17580 19323 17638 19329
rect 17862 19320 17868 19332
rect 17920 19320 17926 19372
rect 19076 19360 19104 19468
rect 20438 19456 20444 19468
rect 20496 19456 20502 19508
rect 24026 19496 24032 19508
rect 22480 19468 24032 19496
rect 19153 19431 19211 19437
rect 19153 19397 19165 19431
rect 19199 19428 19211 19431
rect 22480 19428 22508 19468
rect 24026 19456 24032 19468
rect 24084 19496 24090 19508
rect 24762 19496 24768 19508
rect 24084 19468 24768 19496
rect 24084 19456 24090 19468
rect 24762 19456 24768 19468
rect 24820 19456 24826 19508
rect 27798 19496 27804 19508
rect 27172 19468 27804 19496
rect 19199 19400 22508 19428
rect 22548 19431 22606 19437
rect 19199 19397 19211 19400
rect 19153 19391 19211 19397
rect 22548 19397 22560 19431
rect 22594 19428 22606 19431
rect 23014 19428 23020 19440
rect 22594 19400 23020 19428
rect 22594 19397 22606 19400
rect 22548 19391 22606 19397
rect 23014 19388 23020 19400
rect 23072 19388 23078 19440
rect 24854 19428 24860 19440
rect 24136 19400 24860 19428
rect 19076 19332 19472 19360
rect 19444 19304 19472 19332
rect 20438 19320 20444 19372
rect 20496 19360 20502 19372
rect 22281 19363 22339 19369
rect 22281 19360 22293 19363
rect 20496 19332 22293 19360
rect 20496 19320 20502 19332
rect 22281 19329 22293 19332
rect 22327 19329 22339 19363
rect 23750 19360 23756 19372
rect 22281 19323 22339 19329
rect 23676 19332 23756 19360
rect 16776 19264 16988 19292
rect 19426 19252 19432 19304
rect 19484 19252 19490 19304
rect 16666 19224 16672 19236
rect 16627 19196 16672 19224
rect 16666 19184 16672 19196
rect 16724 19184 16730 19236
rect 23676 19233 23704 19332
rect 23750 19320 23756 19332
rect 23808 19320 23814 19372
rect 24136 19369 24164 19400
rect 24854 19388 24860 19400
rect 24912 19428 24918 19440
rect 25038 19428 25044 19440
rect 24912 19400 25044 19428
rect 24912 19388 24918 19400
rect 25038 19388 25044 19400
rect 25096 19388 25102 19440
rect 26694 19388 26700 19440
rect 26752 19428 26758 19440
rect 27172 19428 27200 19468
rect 27798 19456 27804 19468
rect 27856 19496 27862 19508
rect 28353 19499 28411 19505
rect 28353 19496 28365 19499
rect 27856 19468 28365 19496
rect 27856 19456 27862 19468
rect 28353 19465 28365 19468
rect 28399 19465 28411 19499
rect 30190 19496 30196 19508
rect 30151 19468 30196 19496
rect 28353 19459 28411 19465
rect 30190 19456 30196 19468
rect 30248 19456 30254 19508
rect 32214 19496 32220 19508
rect 32175 19468 32220 19496
rect 32214 19456 32220 19468
rect 32272 19456 32278 19508
rect 33321 19499 33379 19505
rect 33321 19465 33333 19499
rect 33367 19496 33379 19499
rect 34698 19496 34704 19508
rect 33367 19468 34704 19496
rect 33367 19465 33379 19468
rect 33321 19459 33379 19465
rect 34698 19456 34704 19468
rect 34756 19456 34762 19508
rect 34790 19456 34796 19508
rect 34848 19496 34854 19508
rect 35161 19499 35219 19505
rect 35161 19496 35173 19499
rect 34848 19468 35173 19496
rect 34848 19456 34854 19468
rect 35161 19465 35173 19468
rect 35207 19465 35219 19499
rect 35161 19459 35219 19465
rect 26752 19400 27200 19428
rect 26752 19388 26758 19400
rect 27430 19388 27436 19440
rect 27488 19428 27494 19440
rect 29058 19431 29116 19437
rect 29058 19428 29070 19431
rect 27488 19400 29070 19428
rect 27488 19388 27494 19400
rect 29058 19397 29070 19400
rect 29104 19397 29116 19431
rect 34422 19428 34428 19440
rect 29058 19391 29116 19397
rect 33796 19400 34428 19428
rect 24394 19369 24400 19372
rect 24121 19363 24179 19369
rect 24121 19329 24133 19363
rect 24167 19329 24179 19363
rect 24121 19323 24179 19329
rect 24388 19323 24400 19369
rect 24452 19360 24458 19372
rect 25056 19360 25084 19388
rect 26973 19363 27031 19369
rect 26973 19360 26985 19363
rect 24452 19332 24488 19360
rect 25056 19332 26985 19360
rect 24394 19320 24400 19323
rect 24452 19320 24458 19332
rect 26973 19329 26985 19332
rect 27019 19329 27031 19363
rect 26973 19323 27031 19329
rect 27062 19320 27068 19372
rect 27120 19360 27126 19372
rect 27229 19363 27287 19369
rect 27229 19360 27241 19363
rect 27120 19332 27241 19360
rect 27120 19320 27126 19332
rect 27229 19329 27241 19332
rect 27275 19329 27287 19363
rect 28810 19360 28816 19372
rect 28771 19332 28816 19360
rect 27229 19323 27287 19329
rect 28810 19320 28816 19332
rect 28868 19320 28874 19372
rect 30834 19320 30840 19372
rect 30892 19360 30898 19372
rect 30929 19363 30987 19369
rect 30929 19360 30941 19363
rect 30892 19332 30941 19360
rect 30892 19320 30898 19332
rect 30929 19329 30941 19332
rect 30975 19329 30987 19363
rect 32398 19360 32404 19372
rect 32359 19332 32404 19360
rect 30929 19323 30987 19329
rect 32398 19320 32404 19332
rect 32456 19320 32462 19372
rect 33134 19360 33140 19372
rect 33095 19332 33140 19360
rect 33134 19320 33140 19332
rect 33192 19320 33198 19372
rect 33594 19320 33600 19372
rect 33652 19360 33658 19372
rect 33796 19369 33824 19400
rect 34422 19388 34428 19400
rect 34480 19388 34486 19440
rect 33781 19363 33839 19369
rect 33781 19360 33793 19363
rect 33652 19332 33793 19360
rect 33652 19320 33658 19332
rect 33781 19329 33793 19332
rect 33827 19329 33839 19363
rect 33781 19323 33839 19329
rect 34048 19363 34106 19369
rect 34048 19329 34060 19363
rect 34094 19360 34106 19363
rect 34330 19360 34336 19372
rect 34094 19332 34336 19360
rect 34094 19329 34106 19332
rect 34048 19323 34106 19329
rect 34330 19320 34336 19332
rect 34388 19320 34394 19372
rect 37553 19363 37611 19369
rect 37553 19329 37565 19363
rect 37599 19360 37611 19363
rect 37642 19360 37648 19372
rect 37599 19332 37648 19360
rect 37599 19329 37611 19332
rect 37553 19323 37611 19329
rect 37642 19320 37648 19332
rect 37700 19320 37706 19372
rect 32950 19292 32956 19304
rect 32911 19264 32956 19292
rect 32950 19252 32956 19264
rect 33008 19252 33014 19304
rect 37274 19292 37280 19304
rect 37235 19264 37280 19292
rect 37274 19252 37280 19264
rect 37332 19252 37338 19304
rect 23661 19227 23719 19233
rect 23661 19193 23673 19227
rect 23707 19193 23719 19227
rect 23661 19187 23719 19193
rect 4798 19156 4804 19168
rect 4759 19128 4804 19156
rect 4798 19116 4804 19128
rect 4856 19116 4862 19168
rect 7742 19156 7748 19168
rect 7703 19128 7748 19156
rect 7742 19116 7748 19128
rect 7800 19116 7806 19168
rect 10965 19159 11023 19165
rect 10965 19125 10977 19159
rect 11011 19156 11023 19159
rect 11146 19156 11152 19168
rect 11011 19128 11152 19156
rect 11011 19125 11023 19128
rect 10965 19119 11023 19125
rect 11146 19116 11152 19128
rect 11204 19116 11210 19168
rect 15194 19116 15200 19168
rect 15252 19156 15258 19168
rect 16025 19159 16083 19165
rect 16025 19156 16037 19159
rect 15252 19128 16037 19156
rect 15252 19116 15258 19128
rect 16025 19125 16037 19128
rect 16071 19125 16083 19159
rect 16025 19119 16083 19125
rect 24302 19116 24308 19168
rect 24360 19156 24366 19168
rect 25501 19159 25559 19165
rect 25501 19156 25513 19159
rect 24360 19128 25513 19156
rect 24360 19116 24366 19128
rect 25501 19125 25513 19128
rect 25547 19125 25559 19159
rect 30742 19156 30748 19168
rect 30703 19128 30748 19156
rect 25501 19119 25559 19125
rect 30742 19116 30748 19128
rect 30800 19116 30806 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 3786 18912 3792 18964
rect 3844 18952 3850 18964
rect 5445 18955 5503 18961
rect 5445 18952 5457 18955
rect 3844 18924 5457 18952
rect 3844 18912 3850 18924
rect 5445 18921 5457 18924
rect 5491 18952 5503 18955
rect 5534 18952 5540 18964
rect 5491 18924 5540 18952
rect 5491 18921 5503 18924
rect 5445 18915 5503 18921
rect 5534 18912 5540 18924
rect 5592 18912 5598 18964
rect 6641 18955 6699 18961
rect 6641 18921 6653 18955
rect 6687 18952 6699 18955
rect 7742 18952 7748 18964
rect 6687 18924 7748 18952
rect 6687 18921 6699 18924
rect 6641 18915 6699 18921
rect 7742 18912 7748 18924
rect 7800 18912 7806 18964
rect 8113 18955 8171 18961
rect 8113 18921 8125 18955
rect 8159 18952 8171 18955
rect 8662 18952 8668 18964
rect 8159 18924 8668 18952
rect 8159 18921 8171 18924
rect 8113 18915 8171 18921
rect 8662 18912 8668 18924
rect 8720 18912 8726 18964
rect 10321 18955 10379 18961
rect 10321 18921 10333 18955
rect 10367 18952 10379 18955
rect 11054 18952 11060 18964
rect 10367 18924 11060 18952
rect 10367 18921 10379 18924
rect 10321 18915 10379 18921
rect 11054 18912 11060 18924
rect 11112 18912 11118 18964
rect 17586 18952 17592 18964
rect 15672 18924 17592 18952
rect 5810 18844 5816 18896
rect 5868 18884 5874 18896
rect 6825 18887 6883 18893
rect 6825 18884 6837 18887
rect 5868 18856 6837 18884
rect 5868 18844 5874 18856
rect 6825 18853 6837 18856
rect 6871 18853 6883 18887
rect 15562 18884 15568 18896
rect 6825 18847 6883 18853
rect 13280 18856 15568 18884
rect 8386 18816 8392 18828
rect 4172 18788 8392 18816
rect 4172 18757 4200 18788
rect 8386 18776 8392 18788
rect 8444 18816 8450 18828
rect 9214 18816 9220 18828
rect 8444 18788 9220 18816
rect 8444 18776 8450 18788
rect 9214 18776 9220 18788
rect 9272 18776 9278 18828
rect 12618 18816 12624 18828
rect 10704 18788 12624 18816
rect 4157 18751 4215 18757
rect 4157 18717 4169 18751
rect 4203 18717 4215 18751
rect 8294 18748 8300 18760
rect 8255 18720 8300 18748
rect 4157 18711 4215 18717
rect 8294 18708 8300 18720
rect 8352 18708 8358 18760
rect 10502 18708 10508 18760
rect 10560 18748 10566 18760
rect 10704 18757 10732 18788
rect 10597 18751 10655 18757
rect 10597 18748 10609 18751
rect 10560 18720 10609 18748
rect 10560 18708 10566 18720
rect 10597 18717 10609 18720
rect 10643 18717 10655 18751
rect 10597 18711 10655 18717
rect 10689 18751 10747 18757
rect 10689 18717 10701 18751
rect 10735 18717 10747 18751
rect 10689 18711 10747 18717
rect 10781 18751 10839 18757
rect 10781 18717 10793 18751
rect 10827 18717 10839 18751
rect 10781 18711 10839 18717
rect 10965 18751 11023 18757
rect 10965 18717 10977 18751
rect 11011 18717 11023 18751
rect 10965 18711 11023 18717
rect 6454 18680 6460 18692
rect 6415 18652 6460 18680
rect 6454 18640 6460 18652
rect 6512 18640 6518 18692
rect 5350 18572 5356 18624
rect 5408 18612 5414 18624
rect 6657 18615 6715 18621
rect 6657 18612 6669 18615
rect 5408 18584 6669 18612
rect 5408 18572 5414 18584
rect 6657 18581 6669 18584
rect 6703 18581 6715 18615
rect 10796 18612 10824 18711
rect 10980 18680 11008 18711
rect 11054 18708 11060 18760
rect 11112 18748 11118 18760
rect 11808 18757 11836 18788
rect 12618 18776 12624 18788
rect 12676 18776 12682 18828
rect 11701 18751 11759 18757
rect 11701 18748 11713 18751
rect 11112 18720 11713 18748
rect 11112 18708 11118 18720
rect 11701 18717 11713 18720
rect 11747 18717 11759 18751
rect 11701 18711 11759 18717
rect 11793 18751 11851 18757
rect 11793 18717 11805 18751
rect 11839 18717 11851 18751
rect 11793 18711 11851 18717
rect 11885 18751 11943 18757
rect 11885 18717 11897 18751
rect 11931 18717 11943 18751
rect 12066 18748 12072 18760
rect 12027 18720 12072 18748
rect 11885 18711 11943 18717
rect 11900 18680 11928 18711
rect 12066 18708 12072 18720
rect 12124 18708 12130 18760
rect 13170 18748 13176 18760
rect 13131 18720 13176 18748
rect 13170 18708 13176 18720
rect 13228 18708 13234 18760
rect 13280 18757 13308 18856
rect 15562 18844 15568 18856
rect 15620 18844 15626 18896
rect 13814 18816 13820 18828
rect 13372 18788 13820 18816
rect 13372 18757 13400 18788
rect 13814 18776 13820 18788
rect 13872 18776 13878 18828
rect 13998 18776 14004 18828
rect 14056 18816 14062 18828
rect 14369 18819 14427 18825
rect 14369 18816 14381 18819
rect 14056 18788 14381 18816
rect 14056 18776 14062 18788
rect 14369 18785 14381 18788
rect 14415 18785 14427 18819
rect 15672 18816 15700 18924
rect 17586 18912 17592 18924
rect 17644 18952 17650 18964
rect 17644 18924 20852 18952
rect 17644 18912 17650 18924
rect 15746 18844 15752 18896
rect 15804 18884 15810 18896
rect 15804 18856 15884 18884
rect 15804 18844 15810 18856
rect 14369 18779 14427 18785
rect 15120 18788 15700 18816
rect 13265 18751 13323 18757
rect 13265 18717 13277 18751
rect 13311 18717 13323 18751
rect 13265 18711 13323 18717
rect 13357 18751 13415 18757
rect 13357 18717 13369 18751
rect 13403 18717 13415 18751
rect 13357 18711 13415 18717
rect 13541 18751 13599 18757
rect 13541 18717 13553 18751
rect 13587 18748 13599 18751
rect 14093 18751 14151 18757
rect 13587 18720 14044 18748
rect 13587 18717 13599 18720
rect 13541 18711 13599 18717
rect 14016 18692 14044 18720
rect 14093 18717 14105 18751
rect 14139 18748 14151 18751
rect 15120 18748 15148 18788
rect 15746 18748 15752 18760
rect 14139 18720 15148 18748
rect 15707 18720 15752 18748
rect 14139 18717 14151 18720
rect 14093 18711 14151 18717
rect 15746 18708 15752 18720
rect 15804 18708 15810 18760
rect 15856 18757 15884 18856
rect 19242 18844 19248 18896
rect 19300 18884 19306 18896
rect 20824 18884 20852 18924
rect 20898 18912 20904 18964
rect 20956 18952 20962 18964
rect 23201 18955 23259 18961
rect 23201 18952 23213 18955
rect 20956 18924 23213 18952
rect 20956 18912 20962 18924
rect 23201 18921 23213 18924
rect 23247 18921 23259 18955
rect 24394 18952 24400 18964
rect 24355 18924 24400 18952
rect 23201 18915 23259 18921
rect 24394 18912 24400 18924
rect 24452 18912 24458 18964
rect 26513 18955 26571 18961
rect 26513 18921 26525 18955
rect 26559 18952 26571 18955
rect 27062 18952 27068 18964
rect 26559 18924 27068 18952
rect 26559 18921 26571 18924
rect 26513 18915 26571 18921
rect 27062 18912 27068 18924
rect 27120 18912 27126 18964
rect 27890 18912 27896 18964
rect 27948 18952 27954 18964
rect 27985 18955 28043 18961
rect 27985 18952 27997 18955
rect 27948 18924 27997 18952
rect 27948 18912 27954 18924
rect 27985 18921 27997 18924
rect 28031 18921 28043 18955
rect 27985 18915 28043 18921
rect 34057 18955 34115 18961
rect 34057 18921 34069 18955
rect 34103 18952 34115 18955
rect 34514 18952 34520 18964
rect 34103 18924 34520 18952
rect 34103 18921 34115 18924
rect 34057 18915 34115 18921
rect 34514 18912 34520 18924
rect 34572 18912 34578 18964
rect 21634 18884 21640 18896
rect 19300 18856 19840 18884
rect 20824 18856 21640 18884
rect 19300 18844 19306 18856
rect 16574 18816 16580 18828
rect 16040 18788 16580 18816
rect 15841 18751 15899 18757
rect 15841 18717 15853 18751
rect 15887 18717 15899 18751
rect 15841 18711 15899 18717
rect 15933 18751 15991 18757
rect 15933 18717 15945 18751
rect 15979 18748 15991 18751
rect 16040 18748 16068 18788
rect 16574 18776 16580 18788
rect 16632 18776 16638 18828
rect 19334 18816 19340 18828
rect 16684 18788 17264 18816
rect 15979 18720 16068 18748
rect 16117 18751 16175 18757
rect 15979 18717 15991 18720
rect 15933 18711 15991 18717
rect 16117 18717 16129 18751
rect 16163 18748 16175 18751
rect 16206 18748 16212 18760
rect 16163 18720 16212 18748
rect 16163 18717 16175 18720
rect 16117 18711 16175 18717
rect 16206 18708 16212 18720
rect 16264 18708 16270 18760
rect 16684 18748 16712 18788
rect 16850 18748 16856 18760
rect 16316 18720 16712 18748
rect 16811 18720 16856 18748
rect 11974 18680 11980 18692
rect 10980 18652 11980 18680
rect 11974 18640 11980 18652
rect 12032 18640 12038 18692
rect 13998 18640 14004 18692
rect 14056 18680 14062 18692
rect 15010 18680 15016 18692
rect 14056 18652 15016 18680
rect 14056 18640 14062 18652
rect 15010 18640 15016 18652
rect 15068 18680 15074 18692
rect 16316 18680 16344 18720
rect 16850 18708 16856 18720
rect 16908 18708 16914 18760
rect 16945 18751 17003 18757
rect 16945 18717 16957 18751
rect 16991 18717 17003 18751
rect 16945 18711 17003 18717
rect 15068 18652 16344 18680
rect 15068 18640 15074 18652
rect 10962 18612 10968 18624
rect 10796 18584 10968 18612
rect 6657 18575 6715 18581
rect 10962 18572 10968 18584
rect 11020 18572 11026 18624
rect 11425 18615 11483 18621
rect 11425 18581 11437 18615
rect 11471 18612 11483 18615
rect 12250 18612 12256 18624
rect 11471 18584 12256 18612
rect 11471 18581 11483 18584
rect 11425 18575 11483 18581
rect 12250 18572 12256 18584
rect 12308 18572 12314 18624
rect 12894 18612 12900 18624
rect 12855 18584 12900 18612
rect 12894 18572 12900 18584
rect 12952 18572 12958 18624
rect 15473 18615 15531 18621
rect 15473 18581 15485 18615
rect 15519 18612 15531 18615
rect 16298 18612 16304 18624
rect 15519 18584 16304 18612
rect 15519 18581 15531 18584
rect 15473 18575 15531 18581
rect 16298 18572 16304 18584
rect 16356 18572 16362 18624
rect 16574 18612 16580 18624
rect 16535 18584 16580 18612
rect 16574 18572 16580 18584
rect 16632 18572 16638 18624
rect 16960 18612 16988 18711
rect 17034 18708 17040 18760
rect 17092 18748 17098 18760
rect 17236 18757 17264 18788
rect 18432 18788 19340 18816
rect 17221 18751 17279 18757
rect 17092 18720 17137 18748
rect 17092 18708 17098 18720
rect 17221 18717 17233 18751
rect 17267 18717 17279 18751
rect 18322 18748 18328 18760
rect 18283 18720 18328 18748
rect 17221 18711 17279 18717
rect 18322 18708 18328 18720
rect 18380 18708 18386 18760
rect 18432 18757 18460 18788
rect 19334 18776 19340 18788
rect 19392 18776 19398 18828
rect 19812 18825 19840 18856
rect 21634 18844 21640 18856
rect 21692 18884 21698 18896
rect 22094 18884 22100 18896
rect 21692 18856 22100 18884
rect 21692 18844 21698 18856
rect 22094 18844 22100 18856
rect 22152 18884 22158 18896
rect 23106 18884 23112 18896
rect 22152 18856 23112 18884
rect 22152 18844 22158 18856
rect 23106 18844 23112 18856
rect 23164 18844 23170 18896
rect 27338 18884 27344 18896
rect 26896 18856 27344 18884
rect 19797 18819 19855 18825
rect 19797 18785 19809 18819
rect 19843 18785 19855 18819
rect 22557 18819 22615 18825
rect 22557 18816 22569 18819
rect 19797 18779 19855 18785
rect 22112 18788 22569 18816
rect 18417 18751 18475 18757
rect 18417 18717 18429 18751
rect 18463 18717 18475 18751
rect 18417 18711 18475 18717
rect 18509 18751 18567 18757
rect 18509 18717 18521 18751
rect 18555 18748 18567 18751
rect 18598 18748 18604 18760
rect 18555 18720 18604 18748
rect 18555 18717 18567 18720
rect 18509 18711 18567 18717
rect 18598 18708 18604 18720
rect 18656 18708 18662 18760
rect 18690 18708 18696 18760
rect 18748 18748 18754 18760
rect 20073 18751 20131 18757
rect 18748 18720 18793 18748
rect 18748 18708 18754 18720
rect 20073 18717 20085 18751
rect 20119 18748 20131 18751
rect 21315 18751 21373 18757
rect 21441 18754 21447 18760
rect 21315 18748 21327 18751
rect 20119 18720 21327 18748
rect 20119 18717 20131 18720
rect 20073 18711 20131 18717
rect 21315 18717 21327 18720
rect 21361 18717 21373 18751
rect 21315 18711 21373 18717
rect 21434 18748 21447 18754
rect 21434 18714 21446 18748
rect 18340 18680 18368 18708
rect 19978 18680 19984 18692
rect 18340 18652 19984 18680
rect 19978 18640 19984 18652
rect 20036 18680 20042 18692
rect 20088 18680 20116 18711
rect 21434 18708 21447 18714
rect 21499 18708 21505 18760
rect 21545 18751 21603 18757
rect 21545 18717 21557 18751
rect 21591 18717 21603 18751
rect 21545 18711 21603 18717
rect 21741 18751 21799 18757
rect 21741 18717 21753 18751
rect 21787 18748 21799 18751
rect 22002 18748 22008 18760
rect 21787 18720 22008 18748
rect 21787 18717 21799 18720
rect 21741 18711 21799 18717
rect 20036 18652 20116 18680
rect 20036 18640 20042 18652
rect 20346 18640 20352 18692
rect 20404 18680 20410 18692
rect 21560 18680 21588 18711
rect 22002 18708 22008 18720
rect 22060 18708 22066 18760
rect 20404 18652 21312 18680
rect 21560 18652 21680 18680
rect 20404 18640 20410 18652
rect 17218 18612 17224 18624
rect 16960 18584 17224 18612
rect 17218 18572 17224 18584
rect 17276 18572 17282 18624
rect 18049 18615 18107 18621
rect 18049 18581 18061 18615
rect 18095 18612 18107 18615
rect 19058 18612 19064 18624
rect 18095 18584 19064 18612
rect 18095 18581 18107 18584
rect 18049 18575 18107 18581
rect 19058 18572 19064 18584
rect 19116 18572 19122 18624
rect 21085 18615 21143 18621
rect 21085 18581 21097 18615
rect 21131 18612 21143 18615
rect 21174 18612 21180 18624
rect 21131 18584 21180 18612
rect 21131 18581 21143 18584
rect 21085 18575 21143 18581
rect 21174 18572 21180 18584
rect 21232 18572 21238 18624
rect 21284 18612 21312 18652
rect 21652 18612 21680 18652
rect 22112 18612 22140 18788
rect 22557 18785 22569 18788
rect 22603 18785 22615 18819
rect 22557 18779 22615 18785
rect 23566 18776 23572 18828
rect 23624 18816 23630 18828
rect 26896 18816 26924 18856
rect 27338 18844 27344 18856
rect 27396 18844 27402 18896
rect 28166 18816 28172 18828
rect 23624 18788 26924 18816
rect 23624 18776 23630 18788
rect 22370 18748 22376 18760
rect 22331 18720 22376 18748
rect 22370 18708 22376 18720
rect 22428 18708 22434 18760
rect 23290 18708 23296 18760
rect 23348 18748 23354 18760
rect 24780 18757 24808 18788
rect 24673 18751 24731 18757
rect 24673 18748 24685 18751
rect 23348 18720 24685 18748
rect 23348 18708 23354 18720
rect 22189 18683 22247 18689
rect 22189 18649 22201 18683
rect 22235 18649 22247 18683
rect 22189 18643 22247 18649
rect 23109 18683 23167 18689
rect 23109 18649 23121 18683
rect 23155 18680 23167 18683
rect 23198 18680 23204 18692
rect 23155 18652 23204 18680
rect 23155 18649 23167 18652
rect 23109 18643 23167 18649
rect 21284 18584 22140 18612
rect 22204 18612 22232 18643
rect 23198 18640 23204 18652
rect 23256 18640 23262 18692
rect 23382 18612 23388 18624
rect 22204 18584 23388 18612
rect 23382 18572 23388 18584
rect 23440 18572 23446 18624
rect 24412 18612 24440 18720
rect 24673 18717 24685 18720
rect 24719 18717 24731 18751
rect 24673 18711 24731 18717
rect 24765 18751 24823 18757
rect 24765 18717 24777 18751
rect 24811 18717 24823 18751
rect 24765 18711 24823 18717
rect 24857 18751 24915 18757
rect 24857 18717 24869 18751
rect 24903 18717 24915 18751
rect 24857 18711 24915 18717
rect 25041 18751 25099 18757
rect 25041 18717 25053 18751
rect 25087 18748 25099 18751
rect 25222 18748 25228 18760
rect 25087 18720 25228 18748
rect 25087 18717 25099 18720
rect 25041 18711 25099 18717
rect 24486 18640 24492 18692
rect 24544 18680 24550 18692
rect 24872 18680 24900 18711
rect 25222 18708 25228 18720
rect 25280 18708 25286 18760
rect 26602 18708 26608 18760
rect 26660 18748 26666 18760
rect 26896 18757 26924 18788
rect 27172 18788 28172 18816
rect 26789 18751 26847 18757
rect 26789 18748 26801 18751
rect 26660 18720 26801 18748
rect 26660 18708 26666 18720
rect 26789 18717 26801 18720
rect 26835 18717 26847 18751
rect 26789 18711 26847 18717
rect 26881 18751 26939 18757
rect 26881 18717 26893 18751
rect 26927 18717 26939 18751
rect 26881 18711 26939 18717
rect 26970 18708 26976 18760
rect 27028 18748 27034 18760
rect 27172 18757 27200 18788
rect 28166 18776 28172 18788
rect 28224 18776 28230 18828
rect 32585 18819 32643 18825
rect 32585 18785 32597 18819
rect 32631 18816 32643 18819
rect 32950 18816 32956 18828
rect 32631 18788 32956 18816
rect 32631 18785 32643 18788
rect 32585 18779 32643 18785
rect 32950 18776 32956 18788
rect 33008 18776 33014 18828
rect 34698 18816 34704 18828
rect 34659 18788 34704 18816
rect 34698 18776 34704 18788
rect 34756 18776 34762 18828
rect 27157 18751 27215 18757
rect 27028 18720 27073 18748
rect 27028 18708 27034 18720
rect 27157 18717 27169 18751
rect 27203 18717 27215 18751
rect 27157 18711 27215 18717
rect 24544 18652 24900 18680
rect 25240 18680 25268 18708
rect 27172 18680 27200 18711
rect 27246 18708 27252 18760
rect 27304 18748 27310 18760
rect 27617 18751 27675 18757
rect 27617 18748 27629 18751
rect 27304 18720 27629 18748
rect 27304 18708 27310 18720
rect 27617 18717 27629 18720
rect 27663 18717 27675 18751
rect 27617 18711 27675 18717
rect 27801 18751 27859 18757
rect 27801 18717 27813 18751
rect 27847 18748 27859 18751
rect 28074 18748 28080 18760
rect 27847 18720 28080 18748
rect 27847 18717 27859 18720
rect 27801 18711 27859 18717
rect 28074 18708 28080 18720
rect 28132 18708 28138 18760
rect 30650 18748 30656 18760
rect 30611 18720 30656 18748
rect 30650 18708 30656 18720
rect 30708 18708 30714 18760
rect 30742 18708 30748 18760
rect 30800 18748 30806 18760
rect 30909 18751 30967 18757
rect 30909 18748 30921 18751
rect 30800 18720 30921 18748
rect 30800 18708 30806 18720
rect 30909 18717 30921 18720
rect 30955 18717 30967 18751
rect 32766 18748 32772 18760
rect 32727 18720 32772 18748
rect 30909 18711 30967 18717
rect 32766 18708 32772 18720
rect 32824 18708 32830 18760
rect 33134 18708 33140 18760
rect 33192 18748 33198 18760
rect 33873 18751 33931 18757
rect 33873 18748 33885 18751
rect 33192 18720 33885 18748
rect 33192 18708 33198 18720
rect 33873 18717 33885 18720
rect 33919 18717 33931 18751
rect 34974 18748 34980 18760
rect 34935 18720 34980 18748
rect 33873 18711 33931 18717
rect 34974 18708 34980 18720
rect 35032 18708 35038 18760
rect 33686 18680 33692 18692
rect 25240 18652 27200 18680
rect 33647 18652 33692 18680
rect 24544 18640 24550 18652
rect 33686 18640 33692 18652
rect 33744 18640 33750 18692
rect 25222 18612 25228 18624
rect 24412 18584 25228 18612
rect 25222 18572 25228 18584
rect 25280 18572 25286 18624
rect 30926 18572 30932 18624
rect 30984 18612 30990 18624
rect 32033 18615 32091 18621
rect 32033 18612 32045 18615
rect 30984 18584 32045 18612
rect 30984 18572 30990 18584
rect 32033 18581 32045 18584
rect 32079 18581 32091 18615
rect 32033 18575 32091 18581
rect 32953 18615 33011 18621
rect 32953 18581 32965 18615
rect 32999 18612 33011 18615
rect 33042 18612 33048 18624
rect 32999 18584 33048 18612
rect 32999 18581 33011 18584
rect 32953 18575 33011 18581
rect 33042 18572 33048 18584
rect 33100 18572 33106 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 6914 18368 6920 18420
rect 6972 18408 6978 18420
rect 7929 18411 7987 18417
rect 7929 18408 7941 18411
rect 6972 18380 7941 18408
rect 6972 18368 6978 18380
rect 7929 18377 7941 18380
rect 7975 18377 7987 18411
rect 7929 18371 7987 18377
rect 10778 18368 10784 18420
rect 10836 18408 10842 18420
rect 10965 18411 11023 18417
rect 10965 18408 10977 18411
rect 10836 18380 10977 18408
rect 10836 18368 10842 18380
rect 10965 18377 10977 18380
rect 11011 18377 11023 18411
rect 10965 18371 11023 18377
rect 11974 18368 11980 18420
rect 12032 18408 12038 18420
rect 12069 18411 12127 18417
rect 12069 18408 12081 18411
rect 12032 18380 12081 18408
rect 12032 18368 12038 18380
rect 12069 18377 12081 18380
rect 12115 18377 12127 18411
rect 12069 18371 12127 18377
rect 14642 18368 14648 18420
rect 14700 18368 14706 18420
rect 14918 18368 14924 18420
rect 14976 18408 14982 18420
rect 14976 18380 16436 18408
rect 14976 18368 14982 18380
rect 11885 18343 11943 18349
rect 11885 18309 11897 18343
rect 11931 18340 11943 18343
rect 12342 18340 12348 18352
rect 11931 18312 12348 18340
rect 11931 18309 11943 18312
rect 11885 18303 11943 18309
rect 12342 18300 12348 18312
rect 12400 18300 12406 18352
rect 14660 18340 14688 18368
rect 16408 18352 16436 18380
rect 17862 18368 17868 18420
rect 17920 18408 17926 18420
rect 18141 18411 18199 18417
rect 18141 18408 18153 18411
rect 17920 18380 18153 18408
rect 17920 18368 17926 18380
rect 18141 18377 18153 18380
rect 18187 18377 18199 18411
rect 19889 18411 19947 18417
rect 18141 18371 18199 18377
rect 18340 18380 19472 18408
rect 15194 18340 15200 18352
rect 14660 18312 14780 18340
rect 7837 18275 7895 18281
rect 7837 18241 7849 18275
rect 7883 18272 7895 18275
rect 8846 18272 8852 18284
rect 7883 18244 8852 18272
rect 7883 18241 7895 18244
rect 7837 18235 7895 18241
rect 8846 18232 8852 18244
rect 8904 18232 8910 18284
rect 8938 18232 8944 18284
rect 8996 18272 9002 18284
rect 9585 18275 9643 18281
rect 9585 18272 9597 18275
rect 8996 18244 9597 18272
rect 8996 18232 9002 18244
rect 9585 18241 9597 18244
rect 9631 18241 9643 18275
rect 9585 18235 9643 18241
rect 9852 18275 9910 18281
rect 9852 18241 9864 18275
rect 9898 18272 9910 18275
rect 11606 18272 11612 18284
rect 9898 18244 11612 18272
rect 9898 18241 9910 18244
rect 9852 18235 9910 18241
rect 11606 18232 11612 18244
rect 11664 18232 11670 18284
rect 11698 18232 11704 18284
rect 11756 18272 11762 18284
rect 12621 18275 12679 18281
rect 11756 18244 11801 18272
rect 11756 18232 11762 18244
rect 12621 18241 12633 18275
rect 12667 18272 12679 18275
rect 13078 18272 13084 18284
rect 12667 18244 13084 18272
rect 12667 18241 12679 18244
rect 12621 18235 12679 18241
rect 13078 18232 13084 18244
rect 13136 18232 13142 18284
rect 14550 18232 14556 18284
rect 14608 18281 14614 18284
rect 14752 18281 14780 18312
rect 14865 18312 15200 18340
rect 14865 18284 14893 18312
rect 15194 18300 15200 18312
rect 15252 18300 15258 18352
rect 16390 18300 16396 18352
rect 16448 18340 16454 18352
rect 18340 18340 18368 18380
rect 19334 18340 19340 18352
rect 16448 18312 18368 18340
rect 18524 18312 19340 18340
rect 16448 18300 16454 18312
rect 14608 18275 14657 18281
rect 14608 18241 14611 18275
rect 14645 18241 14657 18275
rect 14608 18235 14657 18241
rect 14737 18275 14795 18281
rect 14737 18241 14749 18275
rect 14783 18241 14795 18275
rect 14737 18235 14795 18241
rect 14850 18278 14908 18284
rect 14850 18244 14862 18278
rect 14896 18244 14908 18278
rect 14850 18238 14908 18244
rect 14608 18232 14614 18235
rect 15010 18232 15016 18284
rect 15068 18272 15074 18284
rect 15565 18275 15623 18281
rect 15068 18244 15113 18272
rect 15068 18232 15074 18244
rect 15565 18241 15577 18275
rect 15611 18272 15623 18275
rect 16022 18272 16028 18284
rect 15611 18244 16028 18272
rect 15611 18241 15623 18244
rect 15565 18235 15623 18241
rect 16022 18232 16028 18244
rect 16080 18232 16086 18284
rect 17218 18232 17224 18284
rect 17276 18272 17282 18284
rect 17405 18275 17463 18281
rect 17405 18272 17417 18275
rect 17276 18244 17417 18272
rect 17276 18232 17282 18244
rect 17405 18241 17417 18244
rect 17451 18241 17463 18275
rect 17586 18272 17592 18284
rect 17547 18244 17592 18272
rect 17405 18235 17463 18241
rect 17586 18232 17592 18244
rect 17644 18232 17650 18284
rect 18524 18281 18552 18312
rect 19334 18300 19340 18312
rect 19392 18300 19398 18352
rect 18371 18275 18429 18281
rect 18156 18247 18383 18275
rect 10962 18096 10968 18148
rect 11020 18136 11026 18148
rect 12805 18139 12863 18145
rect 12805 18136 12817 18139
rect 11020 18108 12817 18136
rect 11020 18096 11026 18108
rect 12805 18105 12817 18108
rect 12851 18136 12863 18139
rect 14918 18136 14924 18148
rect 12851 18108 14924 18136
rect 12851 18105 12863 18108
rect 12805 18099 12863 18105
rect 14918 18096 14924 18108
rect 14976 18096 14982 18148
rect 15102 18096 15108 18148
rect 15160 18136 15166 18148
rect 18156 18136 18184 18247
rect 18371 18241 18383 18247
rect 18417 18241 18429 18275
rect 18371 18235 18429 18241
rect 18509 18275 18567 18281
rect 18509 18241 18521 18275
rect 18555 18241 18567 18275
rect 18509 18235 18567 18241
rect 18598 18232 18604 18284
rect 18656 18272 18662 18284
rect 18785 18275 18843 18281
rect 18656 18244 18749 18272
rect 18656 18232 18662 18244
rect 18785 18241 18797 18275
rect 18831 18272 18843 18275
rect 19444 18272 19472 18380
rect 19889 18377 19901 18411
rect 19935 18408 19947 18411
rect 20162 18408 20168 18420
rect 19935 18380 20168 18408
rect 19935 18377 19947 18380
rect 19889 18371 19947 18377
rect 20162 18368 20168 18380
rect 20220 18368 20226 18420
rect 22066 18380 24440 18408
rect 21085 18343 21143 18349
rect 21085 18309 21097 18343
rect 21131 18309 21143 18343
rect 21085 18303 21143 18309
rect 21269 18343 21327 18349
rect 21269 18309 21281 18343
rect 21315 18340 21327 18343
rect 22066 18340 22094 18380
rect 23106 18340 23112 18352
rect 21315 18312 22094 18340
rect 23067 18312 23112 18340
rect 21315 18309 21327 18312
rect 21269 18303 21327 18309
rect 19886 18272 19892 18284
rect 18831 18244 19892 18272
rect 18831 18241 18843 18244
rect 18785 18235 18843 18241
rect 19886 18232 19892 18244
rect 19944 18232 19950 18284
rect 20165 18275 20223 18281
rect 19996 18247 20177 18275
rect 18616 18204 18644 18232
rect 19610 18204 19616 18216
rect 18616 18176 19616 18204
rect 19610 18164 19616 18176
rect 19668 18164 19674 18216
rect 15160 18108 18552 18136
rect 15160 18096 15166 18108
rect 14366 18068 14372 18080
rect 14327 18040 14372 18068
rect 14366 18028 14372 18040
rect 14424 18028 14430 18080
rect 14734 18028 14740 18080
rect 14792 18068 14798 18080
rect 15657 18071 15715 18077
rect 15657 18068 15669 18071
rect 14792 18040 15669 18068
rect 14792 18028 14798 18040
rect 15657 18037 15669 18040
rect 15703 18068 15715 18071
rect 15746 18068 15752 18080
rect 15703 18040 15752 18068
rect 15703 18037 15715 18040
rect 15657 18031 15715 18037
rect 15746 18028 15752 18040
rect 15804 18028 15810 18080
rect 18524 18068 18552 18108
rect 18598 18096 18604 18148
rect 18656 18136 18662 18148
rect 19702 18136 19708 18148
rect 18656 18108 19708 18136
rect 18656 18096 18662 18108
rect 19702 18096 19708 18108
rect 19760 18096 19766 18148
rect 19996 18068 20024 18247
rect 20165 18241 20177 18247
rect 20211 18241 20223 18275
rect 20165 18235 20223 18241
rect 20257 18275 20315 18281
rect 20257 18241 20269 18275
rect 20303 18241 20315 18275
rect 20257 18235 20315 18241
rect 20272 18204 20300 18235
rect 20346 18232 20352 18284
rect 20404 18272 20410 18284
rect 20533 18275 20591 18281
rect 20404 18244 20449 18272
rect 20404 18232 20410 18244
rect 20533 18241 20545 18275
rect 20579 18272 20668 18275
rect 20806 18272 20812 18284
rect 20579 18247 20812 18272
rect 20579 18241 20591 18247
rect 20640 18244 20812 18247
rect 20533 18235 20591 18241
rect 20806 18232 20812 18244
rect 20864 18232 20870 18284
rect 21100 18272 21128 18303
rect 23106 18300 23112 18312
rect 23164 18300 23170 18352
rect 24302 18340 24308 18352
rect 24263 18312 24308 18340
rect 24302 18300 24308 18312
rect 24360 18300 24366 18352
rect 24412 18340 24440 18380
rect 32398 18368 32404 18420
rect 32456 18408 32462 18420
rect 32493 18411 32551 18417
rect 32493 18408 32505 18411
rect 32456 18380 32505 18408
rect 32456 18368 32462 18380
rect 32493 18377 32505 18380
rect 32539 18377 32551 18411
rect 32493 18371 32551 18377
rect 25038 18340 25044 18352
rect 24412 18312 25044 18340
rect 25038 18300 25044 18312
rect 25096 18300 25102 18352
rect 25133 18343 25191 18349
rect 25133 18309 25145 18343
rect 25179 18340 25191 18343
rect 25590 18340 25596 18352
rect 25179 18312 25596 18340
rect 25179 18309 25191 18312
rect 25133 18303 25191 18309
rect 25590 18300 25596 18312
rect 25648 18300 25654 18352
rect 32306 18340 32312 18352
rect 32267 18312 32312 18340
rect 32306 18300 32312 18312
rect 32364 18300 32370 18352
rect 21634 18272 21640 18284
rect 21100 18244 21640 18272
rect 21634 18232 21640 18244
rect 21692 18232 21698 18284
rect 21821 18275 21879 18281
rect 21821 18241 21833 18275
rect 21867 18272 21879 18275
rect 21910 18272 21916 18284
rect 21867 18244 21916 18272
rect 21867 18241 21879 18244
rect 21821 18235 21879 18241
rect 21910 18232 21916 18244
rect 21968 18232 21974 18284
rect 22005 18275 22063 18281
rect 22005 18241 22017 18275
rect 22051 18272 22063 18275
rect 22554 18272 22560 18284
rect 22051 18244 22560 18272
rect 22051 18241 22063 18244
rect 22005 18235 22063 18241
rect 22554 18232 22560 18244
rect 22612 18232 22618 18284
rect 23293 18275 23351 18281
rect 23293 18241 23305 18275
rect 23339 18272 23351 18275
rect 23382 18272 23388 18284
rect 23339 18244 23388 18272
rect 23339 18241 23351 18244
rect 23293 18235 23351 18241
rect 23382 18232 23388 18244
rect 23440 18232 23446 18284
rect 24118 18272 24124 18284
rect 24031 18244 24124 18272
rect 24118 18232 24124 18244
rect 24176 18272 24182 18284
rect 27246 18272 27252 18284
rect 24176 18244 27252 18272
rect 24176 18232 24182 18244
rect 27246 18232 27252 18244
rect 27304 18232 27310 18284
rect 30466 18232 30472 18284
rect 30524 18272 30530 18284
rect 30653 18275 30711 18281
rect 30653 18272 30665 18275
rect 30524 18244 30665 18272
rect 30524 18232 30530 18244
rect 30653 18241 30665 18244
rect 30699 18241 30711 18275
rect 30926 18272 30932 18284
rect 30887 18244 30932 18272
rect 30653 18235 30711 18241
rect 30926 18232 30932 18244
rect 30984 18232 30990 18284
rect 32122 18272 32128 18284
rect 32083 18244 32128 18272
rect 32122 18232 32128 18244
rect 32180 18232 32186 18284
rect 33042 18272 33048 18284
rect 33003 18244 33048 18272
rect 33042 18232 33048 18244
rect 33100 18232 33106 18284
rect 21450 18204 21456 18216
rect 20272 18176 21456 18204
rect 21450 18164 21456 18176
rect 21508 18164 21514 18216
rect 32950 18204 32956 18216
rect 31726 18176 32956 18204
rect 20898 18136 20904 18148
rect 20732 18108 20904 18136
rect 20732 18068 20760 18108
rect 20898 18096 20904 18108
rect 20956 18096 20962 18148
rect 21266 18096 21272 18148
rect 21324 18136 21330 18148
rect 22189 18139 22247 18145
rect 22189 18136 22201 18139
rect 21324 18108 22201 18136
rect 21324 18096 21330 18108
rect 22189 18105 22201 18108
rect 22235 18105 22247 18139
rect 24486 18136 24492 18148
rect 24447 18108 24492 18136
rect 22189 18099 22247 18105
rect 24486 18096 24492 18108
rect 24544 18096 24550 18148
rect 24670 18096 24676 18148
rect 24728 18136 24734 18148
rect 31726 18136 31754 18176
rect 32950 18164 32956 18176
rect 33008 18164 33014 18216
rect 33321 18207 33379 18213
rect 33321 18173 33333 18207
rect 33367 18204 33379 18207
rect 33502 18204 33508 18216
rect 33367 18176 33508 18204
rect 33367 18173 33379 18176
rect 33321 18167 33379 18173
rect 33502 18164 33508 18176
rect 33560 18164 33566 18216
rect 34514 18164 34520 18216
rect 34572 18204 34578 18216
rect 37277 18207 37335 18213
rect 37277 18204 37289 18207
rect 34572 18176 37289 18204
rect 34572 18164 34578 18176
rect 37277 18173 37289 18176
rect 37323 18173 37335 18207
rect 37277 18167 37335 18173
rect 37553 18207 37611 18213
rect 37553 18173 37565 18207
rect 37599 18204 37611 18207
rect 37826 18204 37832 18216
rect 37599 18176 37832 18204
rect 37599 18173 37611 18176
rect 37553 18167 37611 18173
rect 37826 18164 37832 18176
rect 37884 18164 37890 18216
rect 24728 18108 31754 18136
rect 24728 18096 24734 18108
rect 18524 18040 20760 18068
rect 21726 18028 21732 18080
rect 21784 18068 21790 18080
rect 22002 18068 22008 18080
rect 21784 18040 22008 18068
rect 21784 18028 21790 18040
rect 22002 18028 22008 18040
rect 22060 18028 22066 18080
rect 23290 18028 23296 18080
rect 23348 18068 23354 18080
rect 25130 18068 25136 18080
rect 23348 18040 25136 18068
rect 23348 18028 23354 18040
rect 25130 18028 25136 18040
rect 25188 18068 25194 18080
rect 25225 18071 25283 18077
rect 25225 18068 25237 18071
rect 25188 18040 25237 18068
rect 25188 18028 25194 18040
rect 25225 18037 25237 18040
rect 25271 18037 25283 18071
rect 25225 18031 25283 18037
rect 30469 18071 30527 18077
rect 30469 18037 30481 18071
rect 30515 18068 30527 18071
rect 30558 18068 30564 18080
rect 30515 18040 30564 18068
rect 30515 18037 30527 18040
rect 30469 18031 30527 18037
rect 30558 18028 30564 18040
rect 30616 18028 30622 18080
rect 30742 18028 30748 18080
rect 30800 18068 30806 18080
rect 30837 18071 30895 18077
rect 30837 18068 30849 18071
rect 30800 18040 30849 18068
rect 30800 18028 30806 18040
rect 30837 18037 30849 18040
rect 30883 18037 30895 18071
rect 30837 18031 30895 18037
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 8846 17824 8852 17876
rect 8904 17864 8910 17876
rect 9493 17867 9551 17873
rect 9493 17864 9505 17867
rect 8904 17836 9505 17864
rect 8904 17824 8910 17836
rect 9493 17833 9505 17836
rect 9539 17833 9551 17867
rect 11514 17864 11520 17876
rect 9493 17827 9551 17833
rect 11072 17836 11520 17864
rect 5902 17756 5908 17808
rect 5960 17796 5966 17808
rect 6917 17799 6975 17805
rect 6917 17796 6929 17799
rect 5960 17768 6929 17796
rect 5960 17756 5966 17768
rect 6917 17765 6929 17768
rect 6963 17765 6975 17799
rect 6917 17759 6975 17765
rect 9398 17756 9404 17808
rect 9456 17796 9462 17808
rect 11072 17796 11100 17836
rect 11514 17824 11520 17836
rect 11572 17824 11578 17876
rect 11606 17824 11612 17876
rect 11664 17864 11670 17876
rect 11793 17867 11851 17873
rect 11793 17864 11805 17867
rect 11664 17836 11805 17864
rect 11664 17824 11670 17836
rect 11793 17833 11805 17836
rect 11839 17833 11851 17867
rect 11793 17827 11851 17833
rect 13170 17824 13176 17876
rect 13228 17864 13234 17876
rect 14550 17864 14556 17876
rect 13228 17836 14556 17864
rect 13228 17824 13234 17836
rect 14550 17824 14556 17836
rect 14608 17864 14614 17876
rect 15841 17867 15899 17873
rect 15841 17864 15853 17867
rect 14608 17836 15853 17864
rect 14608 17824 14614 17836
rect 15841 17833 15853 17836
rect 15887 17864 15899 17867
rect 16850 17864 16856 17876
rect 15887 17836 16856 17864
rect 15887 17833 15899 17836
rect 15841 17827 15899 17833
rect 16850 17824 16856 17836
rect 16908 17824 16914 17876
rect 19610 17864 19616 17876
rect 19571 17836 19616 17864
rect 19610 17824 19616 17836
rect 19668 17824 19674 17876
rect 20714 17864 20720 17876
rect 19720 17836 20720 17864
rect 9456 17768 11100 17796
rect 9456 17756 9462 17768
rect 11146 17756 11152 17808
rect 11204 17796 11210 17808
rect 15197 17799 15255 17805
rect 11204 17768 12296 17796
rect 11204 17756 11210 17768
rect 11072 17700 12204 17728
rect 5810 17620 5816 17672
rect 5868 17660 5874 17672
rect 6457 17663 6515 17669
rect 6457 17660 6469 17663
rect 5868 17632 6469 17660
rect 5868 17620 5874 17632
rect 6457 17629 6469 17632
rect 6503 17629 6515 17663
rect 7098 17660 7104 17672
rect 7059 17632 7104 17660
rect 6457 17623 6515 17629
rect 7098 17620 7104 17632
rect 7156 17620 7162 17672
rect 10962 17660 10968 17672
rect 10923 17632 10968 17660
rect 10962 17620 10968 17632
rect 11020 17620 11026 17672
rect 11072 17669 11100 17700
rect 11057 17663 11115 17669
rect 11057 17629 11069 17663
rect 11103 17629 11115 17663
rect 11057 17623 11115 17629
rect 11146 17620 11152 17672
rect 11204 17660 11210 17672
rect 11330 17660 11336 17672
rect 11204 17632 11249 17660
rect 11291 17632 11336 17660
rect 11204 17620 11210 17632
rect 11330 17620 11336 17632
rect 11388 17660 11394 17672
rect 11974 17660 11980 17672
rect 11388 17632 11980 17660
rect 11388 17620 11394 17632
rect 11974 17620 11980 17632
rect 12032 17620 12038 17672
rect 12176 17669 12204 17700
rect 12268 17669 12296 17768
rect 15197 17765 15209 17799
rect 15243 17796 15255 17799
rect 15286 17796 15292 17808
rect 15243 17768 15292 17796
rect 15243 17765 15255 17768
rect 15197 17759 15255 17765
rect 15286 17756 15292 17768
rect 15344 17756 15350 17808
rect 12802 17688 12808 17740
rect 12860 17728 12866 17740
rect 12897 17731 12955 17737
rect 12897 17728 12909 17731
rect 12860 17700 12909 17728
rect 12860 17688 12866 17700
rect 12897 17697 12909 17700
rect 12943 17697 12955 17731
rect 12897 17691 12955 17697
rect 13446 17688 13452 17740
rect 13504 17728 13510 17740
rect 19720 17728 19748 17836
rect 20714 17824 20720 17836
rect 20772 17824 20778 17876
rect 22554 17864 22560 17876
rect 22515 17836 22560 17864
rect 22554 17824 22560 17836
rect 22612 17824 22618 17876
rect 23290 17824 23296 17876
rect 23348 17864 23354 17876
rect 30834 17864 30840 17876
rect 23348 17836 28994 17864
rect 30795 17836 30840 17864
rect 23348 17824 23354 17836
rect 20438 17756 20444 17808
rect 20496 17756 20502 17808
rect 13504 17700 19748 17728
rect 20456 17728 20484 17756
rect 21177 17731 21235 17737
rect 21177 17728 21189 17731
rect 20456 17700 21189 17728
rect 13504 17688 13510 17700
rect 21177 17697 21189 17700
rect 21223 17697 21235 17731
rect 22572 17728 22600 17824
rect 23017 17731 23075 17737
rect 23017 17728 23029 17731
rect 22572 17700 23029 17728
rect 21177 17691 21235 17697
rect 23017 17697 23029 17700
rect 23063 17697 23075 17731
rect 24854 17728 24860 17740
rect 24815 17700 24860 17728
rect 23017 17691 23075 17697
rect 24854 17688 24860 17700
rect 24912 17688 24918 17740
rect 28166 17688 28172 17740
rect 28224 17728 28230 17740
rect 28445 17731 28503 17737
rect 28445 17728 28457 17731
rect 28224 17700 28457 17728
rect 28224 17688 28230 17700
rect 28445 17697 28457 17700
rect 28491 17697 28503 17731
rect 28626 17728 28632 17740
rect 28587 17700 28632 17728
rect 28445 17691 28503 17697
rect 28626 17688 28632 17700
rect 28684 17688 28690 17740
rect 28966 17728 28994 17836
rect 30834 17824 30840 17836
rect 30892 17824 30898 17876
rect 33413 17867 33471 17873
rect 33413 17833 33425 17867
rect 33459 17864 33471 17867
rect 34514 17864 34520 17876
rect 33459 17836 34520 17864
rect 33459 17833 33471 17836
rect 33413 17827 33471 17833
rect 34514 17824 34520 17836
rect 34572 17824 34578 17876
rect 31573 17731 31631 17737
rect 31573 17728 31585 17731
rect 28966 17700 31585 17728
rect 31573 17697 31585 17700
rect 31619 17728 31631 17731
rect 32122 17728 32128 17740
rect 31619 17700 32128 17728
rect 31619 17697 31631 17700
rect 31573 17691 31631 17697
rect 32122 17688 32128 17700
rect 32180 17688 32186 17740
rect 32306 17688 32312 17740
rect 32364 17728 32370 17740
rect 32364 17700 33272 17728
rect 32364 17688 32370 17700
rect 12069 17663 12127 17669
rect 12069 17629 12081 17663
rect 12115 17629 12127 17663
rect 12069 17623 12127 17629
rect 12161 17663 12219 17669
rect 12161 17629 12173 17663
rect 12207 17629 12219 17663
rect 12161 17623 12219 17629
rect 12253 17663 12311 17669
rect 12253 17629 12265 17663
rect 12299 17629 12311 17663
rect 12253 17623 12311 17629
rect 12437 17663 12495 17669
rect 12437 17629 12449 17663
rect 12483 17660 12495 17663
rect 12618 17660 12624 17672
rect 12483 17632 12624 17660
rect 12483 17629 12495 17632
rect 12437 17623 12495 17629
rect 9398 17592 9404 17604
rect 9359 17564 9404 17592
rect 9398 17552 9404 17564
rect 9456 17552 9462 17604
rect 12084 17536 12112 17623
rect 12176 17592 12204 17623
rect 12618 17620 12624 17632
rect 12676 17620 12682 17672
rect 13081 17663 13139 17669
rect 13081 17629 13093 17663
rect 13127 17660 13139 17663
rect 13814 17660 13820 17672
rect 13127 17632 13820 17660
rect 13127 17629 13139 17632
rect 13081 17623 13139 17629
rect 13814 17620 13820 17632
rect 13872 17620 13878 17672
rect 15470 17660 15476 17672
rect 13924 17632 15476 17660
rect 13924 17592 13952 17632
rect 15470 17620 15476 17632
rect 15528 17620 15534 17672
rect 16485 17663 16543 17669
rect 16485 17629 16497 17663
rect 16531 17660 16543 17663
rect 17586 17660 17592 17672
rect 16531 17632 17592 17660
rect 16531 17629 16543 17632
rect 16485 17623 16543 17629
rect 17586 17620 17592 17632
rect 17644 17620 17650 17672
rect 19426 17660 19432 17672
rect 19387 17632 19432 17660
rect 19426 17620 19432 17632
rect 19484 17620 19490 17672
rect 20070 17620 20076 17672
rect 20128 17660 20134 17672
rect 20349 17663 20407 17669
rect 20349 17660 20361 17663
rect 20128 17632 20361 17660
rect 20128 17620 20134 17632
rect 20349 17629 20361 17632
rect 20395 17629 20407 17663
rect 20349 17623 20407 17629
rect 20441 17663 20499 17669
rect 20441 17629 20453 17663
rect 20487 17629 20499 17663
rect 20441 17623 20499 17629
rect 20533 17663 20591 17669
rect 20533 17629 20545 17663
rect 20579 17629 20591 17663
rect 20533 17623 20591 17629
rect 15010 17592 15016 17604
rect 12176 17564 13952 17592
rect 14971 17564 15016 17592
rect 15010 17552 15016 17564
rect 15068 17552 15074 17604
rect 15749 17595 15807 17601
rect 15749 17561 15761 17595
rect 15795 17592 15807 17595
rect 16022 17592 16028 17604
rect 15795 17564 16028 17592
rect 15795 17561 15807 17564
rect 15749 17555 15807 17561
rect 16022 17552 16028 17564
rect 16080 17552 16086 17604
rect 17218 17592 17224 17604
rect 17179 17564 17224 17592
rect 17218 17552 17224 17564
rect 17276 17552 17282 17604
rect 19245 17595 19303 17601
rect 19245 17561 19257 17595
rect 19291 17592 19303 17595
rect 19334 17592 19340 17604
rect 19291 17564 19340 17592
rect 19291 17561 19303 17564
rect 19245 17555 19303 17561
rect 19334 17552 19340 17564
rect 19392 17552 19398 17604
rect 6178 17484 6184 17536
rect 6236 17524 6242 17536
rect 6273 17527 6331 17533
rect 6273 17524 6285 17527
rect 6236 17496 6285 17524
rect 6236 17484 6242 17496
rect 6273 17493 6285 17496
rect 6319 17493 6331 17527
rect 6273 17487 6331 17493
rect 9950 17484 9956 17536
rect 10008 17524 10014 17536
rect 10689 17527 10747 17533
rect 10689 17524 10701 17527
rect 10008 17496 10701 17524
rect 10008 17484 10014 17496
rect 10689 17493 10701 17496
rect 10735 17493 10747 17527
rect 10689 17487 10747 17493
rect 12066 17484 12072 17536
rect 12124 17484 12130 17536
rect 13078 17484 13084 17536
rect 13136 17524 13142 17536
rect 13265 17527 13323 17533
rect 13265 17524 13277 17527
rect 13136 17496 13277 17524
rect 13136 17484 13142 17496
rect 13265 17493 13277 17496
rect 13311 17493 13323 17527
rect 13265 17487 13323 17493
rect 16206 17484 16212 17536
rect 16264 17524 16270 17536
rect 16577 17527 16635 17533
rect 16577 17524 16589 17527
rect 16264 17496 16589 17524
rect 16264 17484 16270 17496
rect 16577 17493 16589 17496
rect 16623 17493 16635 17527
rect 16577 17487 16635 17493
rect 17126 17484 17132 17536
rect 17184 17524 17190 17536
rect 17313 17527 17371 17533
rect 17313 17524 17325 17527
rect 17184 17496 17325 17524
rect 17184 17484 17190 17496
rect 17313 17493 17325 17496
rect 17359 17493 17371 17527
rect 17313 17487 17371 17493
rect 20073 17527 20131 17533
rect 20073 17493 20085 17527
rect 20119 17524 20131 17527
rect 20346 17524 20352 17536
rect 20119 17496 20352 17524
rect 20119 17493 20131 17496
rect 20073 17487 20131 17493
rect 20346 17484 20352 17496
rect 20404 17484 20410 17536
rect 20456 17524 20484 17623
rect 20548 17592 20576 17623
rect 20714 17620 20720 17672
rect 20772 17660 20778 17672
rect 21726 17660 21732 17672
rect 20772 17632 21732 17660
rect 20772 17620 20778 17632
rect 21726 17620 21732 17632
rect 21784 17620 21790 17672
rect 23198 17660 23204 17672
rect 23159 17632 23204 17660
rect 23198 17620 23204 17632
rect 23256 17620 23262 17672
rect 28350 17660 28356 17672
rect 28311 17632 28356 17660
rect 28350 17620 28356 17632
rect 28408 17620 28414 17672
rect 29641 17663 29699 17669
rect 29641 17629 29653 17663
rect 29687 17660 29699 17663
rect 30469 17663 30527 17669
rect 30469 17660 30481 17663
rect 29687 17632 30481 17660
rect 29687 17629 29699 17632
rect 29641 17623 29699 17629
rect 30469 17629 30481 17632
rect 30515 17660 30527 17663
rect 31849 17663 31907 17669
rect 30515 17632 30788 17660
rect 30515 17629 30527 17632
rect 30469 17623 30527 17629
rect 21266 17592 21272 17604
rect 20548 17564 21272 17592
rect 21266 17552 21272 17564
rect 21324 17552 21330 17604
rect 21444 17595 21502 17601
rect 21444 17561 21456 17595
rect 21490 17592 21502 17595
rect 22462 17592 22468 17604
rect 21490 17564 22468 17592
rect 21490 17561 21502 17564
rect 21444 17555 21502 17561
rect 22462 17552 22468 17564
rect 22520 17552 22526 17604
rect 25124 17595 25182 17601
rect 25124 17561 25136 17595
rect 25170 17592 25182 17595
rect 26970 17592 26976 17604
rect 25170 17564 26976 17592
rect 25170 17561 25182 17564
rect 25124 17555 25182 17561
rect 26970 17552 26976 17564
rect 27028 17552 27034 17604
rect 29825 17595 29883 17601
rect 29825 17561 29837 17595
rect 29871 17592 29883 17595
rect 29871 17564 30512 17592
rect 29871 17561 29883 17564
rect 29825 17555 29883 17561
rect 30484 17536 30512 17564
rect 30558 17552 30564 17604
rect 30616 17592 30622 17604
rect 30653 17595 30711 17601
rect 30653 17592 30665 17595
rect 30616 17564 30665 17592
rect 30616 17552 30622 17564
rect 30653 17561 30665 17564
rect 30699 17561 30711 17595
rect 30760 17592 30788 17632
rect 31849 17629 31861 17663
rect 31895 17629 31907 17663
rect 31849 17623 31907 17629
rect 31864 17592 31892 17623
rect 32950 17620 32956 17672
rect 33008 17660 33014 17672
rect 33244 17669 33272 17700
rect 33045 17663 33103 17669
rect 33045 17660 33057 17663
rect 33008 17632 33057 17660
rect 33008 17620 33014 17632
rect 33045 17629 33057 17632
rect 33091 17629 33103 17663
rect 33045 17623 33103 17629
rect 33229 17663 33287 17669
rect 33229 17629 33241 17663
rect 33275 17629 33287 17663
rect 33229 17623 33287 17629
rect 34422 17620 34428 17672
rect 34480 17660 34486 17672
rect 34701 17663 34759 17669
rect 34701 17660 34713 17663
rect 34480 17632 34713 17660
rect 34480 17620 34486 17632
rect 34701 17629 34713 17632
rect 34747 17629 34759 17663
rect 34701 17623 34759 17629
rect 33686 17592 33692 17604
rect 30760 17564 33692 17592
rect 30653 17555 30711 17561
rect 33686 17552 33692 17564
rect 33744 17552 33750 17604
rect 34946 17595 35004 17601
rect 34946 17592 34958 17595
rect 33796 17564 34958 17592
rect 21634 17524 21640 17536
rect 20456 17496 21640 17524
rect 21634 17484 21640 17496
rect 21692 17484 21698 17536
rect 22554 17484 22560 17536
rect 22612 17524 22618 17536
rect 23385 17527 23443 17533
rect 23385 17524 23397 17527
rect 22612 17496 23397 17524
rect 22612 17484 22618 17496
rect 23385 17493 23397 17496
rect 23431 17493 23443 17527
rect 23385 17487 23443 17493
rect 26142 17484 26148 17536
rect 26200 17524 26206 17536
rect 26237 17527 26295 17533
rect 26237 17524 26249 17527
rect 26200 17496 26249 17524
rect 26200 17484 26206 17496
rect 26237 17493 26249 17496
rect 26283 17493 26295 17527
rect 26237 17487 26295 17493
rect 28629 17527 28687 17533
rect 28629 17493 28641 17527
rect 28675 17524 28687 17527
rect 28902 17524 28908 17536
rect 28675 17496 28908 17524
rect 28675 17493 28687 17496
rect 28629 17487 28687 17493
rect 28902 17484 28908 17496
rect 28960 17484 28966 17536
rect 29914 17484 29920 17536
rect 29972 17524 29978 17536
rect 30009 17527 30067 17533
rect 30009 17524 30021 17527
rect 29972 17496 30021 17524
rect 29972 17484 29978 17496
rect 30009 17493 30021 17496
rect 30055 17493 30067 17527
rect 30009 17487 30067 17493
rect 30466 17484 30472 17536
rect 30524 17484 30530 17536
rect 33134 17484 33140 17536
rect 33192 17524 33198 17536
rect 33796 17524 33824 17564
rect 34946 17561 34958 17564
rect 34992 17561 35004 17595
rect 34946 17555 35004 17561
rect 36078 17524 36084 17536
rect 33192 17496 33824 17524
rect 36039 17496 36084 17524
rect 33192 17484 33198 17496
rect 36078 17484 36084 17496
rect 36136 17484 36142 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 4062 17280 4068 17332
rect 4120 17320 4126 17332
rect 7193 17323 7251 17329
rect 7193 17320 7205 17323
rect 4120 17292 7205 17320
rect 4120 17280 4126 17292
rect 7193 17289 7205 17292
rect 7239 17289 7251 17323
rect 12526 17320 12532 17332
rect 12487 17292 12532 17320
rect 7193 17283 7251 17289
rect 12526 17280 12532 17292
rect 12584 17280 12590 17332
rect 12986 17280 12992 17332
rect 13044 17320 13050 17332
rect 13446 17320 13452 17332
rect 13044 17292 13452 17320
rect 13044 17280 13050 17292
rect 13446 17280 13452 17292
rect 13504 17280 13510 17332
rect 15010 17280 15016 17332
rect 15068 17280 15074 17332
rect 18371 17323 18429 17329
rect 18371 17289 18383 17323
rect 18417 17320 18429 17323
rect 18690 17320 18696 17332
rect 18417 17292 18696 17320
rect 18417 17289 18429 17292
rect 18371 17283 18429 17289
rect 18690 17280 18696 17292
rect 18748 17280 18754 17332
rect 20070 17320 20076 17332
rect 19698 17292 20076 17320
rect 6086 17212 6092 17264
rect 6144 17252 6150 17264
rect 6549 17255 6607 17261
rect 6549 17252 6561 17255
rect 6144 17224 6561 17252
rect 6144 17212 6150 17224
rect 6549 17221 6561 17224
rect 6595 17221 6607 17255
rect 6549 17215 6607 17221
rect 6733 17255 6791 17261
rect 6733 17221 6745 17255
rect 6779 17252 6791 17255
rect 11701 17255 11759 17261
rect 6779 17224 8064 17252
rect 6779 17221 6791 17224
rect 6733 17215 6791 17221
rect 2952 17187 3010 17193
rect 2952 17153 2964 17187
rect 2998 17184 3010 17187
rect 5442 17184 5448 17196
rect 2998 17156 5448 17184
rect 2998 17153 3010 17156
rect 2952 17147 3010 17153
rect 5442 17144 5448 17156
rect 5500 17144 5506 17196
rect 5813 17187 5871 17193
rect 5813 17153 5825 17187
rect 5859 17153 5871 17187
rect 5813 17147 5871 17153
rect 6365 17187 6423 17193
rect 6365 17153 6377 17187
rect 6411 17184 6423 17187
rect 7006 17184 7012 17196
rect 6411 17156 7012 17184
rect 6411 17153 6423 17156
rect 6365 17147 6423 17153
rect 2682 17116 2688 17128
rect 2643 17088 2688 17116
rect 2682 17076 2688 17088
rect 2740 17076 2746 17128
rect 3694 17076 3700 17128
rect 3752 17116 3758 17128
rect 5828 17116 5856 17147
rect 7006 17144 7012 17156
rect 7064 17144 7070 17196
rect 7374 17184 7380 17196
rect 7335 17156 7380 17184
rect 7374 17144 7380 17156
rect 7432 17144 7438 17196
rect 8036 17193 8064 17224
rect 11701 17221 11713 17255
rect 11747 17252 11759 17255
rect 13078 17252 13084 17264
rect 11747 17224 13084 17252
rect 11747 17221 11759 17224
rect 11701 17215 11759 17221
rect 13078 17212 13084 17224
rect 13136 17212 13142 17264
rect 13173 17255 13231 17261
rect 13173 17221 13185 17255
rect 13219 17252 13231 17255
rect 14369 17255 14427 17261
rect 13219 17224 14228 17252
rect 13219 17221 13231 17224
rect 13173 17215 13231 17221
rect 8021 17187 8079 17193
rect 8021 17153 8033 17187
rect 8067 17153 8079 17187
rect 8021 17147 8079 17153
rect 8665 17187 8723 17193
rect 8665 17153 8677 17187
rect 8711 17184 8723 17187
rect 9306 17184 9312 17196
rect 8711 17156 9312 17184
rect 8711 17153 8723 17156
rect 8665 17147 8723 17153
rect 9306 17144 9312 17156
rect 9364 17144 9370 17196
rect 12345 17187 12403 17193
rect 12345 17153 12357 17187
rect 12391 17184 12403 17187
rect 13188 17184 13216 17215
rect 12391 17156 13216 17184
rect 12391 17153 12403 17156
rect 12345 17147 12403 17153
rect 8110 17116 8116 17128
rect 3752 17088 5764 17116
rect 5828 17088 8116 17116
rect 3752 17076 3758 17088
rect 4614 17008 4620 17060
rect 4672 17048 4678 17060
rect 5629 17051 5687 17057
rect 5629 17048 5641 17051
rect 4672 17020 5641 17048
rect 4672 17008 4678 17020
rect 5629 17017 5641 17020
rect 5675 17017 5687 17051
rect 5736 17048 5764 17088
rect 8110 17076 8116 17088
rect 8168 17076 8174 17128
rect 8846 17076 8852 17128
rect 8904 17116 8910 17128
rect 12360 17116 12388 17147
rect 13814 17144 13820 17196
rect 13872 17184 13878 17196
rect 14200 17193 14228 17224
rect 14369 17221 14381 17255
rect 14415 17252 14427 17255
rect 15028 17252 15056 17280
rect 15746 17252 15752 17264
rect 14415 17224 15752 17252
rect 14415 17221 14427 17224
rect 14369 17215 14427 17221
rect 15746 17212 15752 17224
rect 15804 17212 15810 17264
rect 16022 17212 16028 17264
rect 16080 17252 16086 17264
rect 16080 17224 18644 17252
rect 16080 17212 16086 17224
rect 14093 17187 14151 17193
rect 14093 17184 14105 17187
rect 13872 17156 14105 17184
rect 13872 17144 13878 17156
rect 14093 17153 14105 17156
rect 14139 17153 14151 17187
rect 14093 17147 14151 17153
rect 14185 17187 14243 17193
rect 14185 17153 14197 17187
rect 14231 17153 14243 17187
rect 14185 17147 14243 17153
rect 8904 17088 12388 17116
rect 14108 17116 14136 17147
rect 14274 17144 14280 17196
rect 14332 17184 14338 17196
rect 15010 17184 15016 17196
rect 14332 17156 15016 17184
rect 14332 17144 14338 17156
rect 15010 17144 15016 17156
rect 15068 17184 15074 17196
rect 15105 17187 15163 17193
rect 15105 17184 15117 17187
rect 15068 17156 15117 17184
rect 15068 17144 15074 17156
rect 15105 17153 15117 17156
rect 15151 17153 15163 17187
rect 15105 17147 15163 17153
rect 15197 17187 15255 17193
rect 15197 17153 15209 17187
rect 15243 17153 15255 17187
rect 15378 17184 15384 17196
rect 15339 17156 15384 17184
rect 15197 17147 15255 17153
rect 14550 17116 14556 17128
rect 14108 17088 14556 17116
rect 8904 17076 8910 17088
rect 14550 17076 14556 17088
rect 14608 17076 14614 17128
rect 15212 17116 15240 17147
rect 15378 17144 15384 17156
rect 15436 17144 15442 17196
rect 15470 17144 15476 17196
rect 15528 17184 15534 17196
rect 15930 17184 15936 17196
rect 15528 17156 15573 17184
rect 15891 17156 15936 17184
rect 15528 17144 15534 17156
rect 15930 17144 15936 17156
rect 15988 17144 15994 17196
rect 17144 17193 17172 17224
rect 17129 17187 17187 17193
rect 17129 17153 17141 17187
rect 17175 17153 17187 17187
rect 17129 17147 17187 17153
rect 17313 17187 17371 17193
rect 17313 17153 17325 17187
rect 17359 17184 17371 17187
rect 17862 17184 17868 17196
rect 17359 17156 17868 17184
rect 17359 17153 17371 17156
rect 17313 17147 17371 17153
rect 17862 17144 17868 17156
rect 17920 17144 17926 17196
rect 18616 17128 18644 17224
rect 18708 17184 18736 17280
rect 19518 17184 19524 17196
rect 18708 17156 19524 17184
rect 19518 17144 19524 17156
rect 19576 17144 19582 17196
rect 19698 17193 19726 17292
rect 20070 17280 20076 17292
rect 20128 17280 20134 17332
rect 20806 17280 20812 17332
rect 20864 17320 20870 17332
rect 20864 17292 21220 17320
rect 20864 17280 20870 17292
rect 20530 17252 20536 17264
rect 19812 17224 20536 17252
rect 19812 17193 19840 17224
rect 20530 17212 20536 17224
rect 20588 17252 20594 17264
rect 20588 17224 20944 17252
rect 20588 17212 20594 17224
rect 19698 17187 19763 17193
rect 19698 17154 19717 17187
rect 19705 17153 19717 17154
rect 19751 17153 19763 17187
rect 19705 17147 19763 17153
rect 19797 17187 19855 17193
rect 19797 17153 19809 17187
rect 19843 17153 19855 17187
rect 19797 17147 19855 17153
rect 19889 17187 19947 17193
rect 19889 17153 19901 17187
rect 19935 17153 19947 17187
rect 19889 17147 19947 17153
rect 20067 17187 20125 17193
rect 20162 17187 20168 17196
rect 20067 17153 20079 17187
rect 20113 17159 20168 17187
rect 20113 17153 20125 17159
rect 20067 17147 20125 17153
rect 15562 17116 15568 17128
rect 15212 17088 15568 17116
rect 15562 17076 15568 17088
rect 15620 17076 15626 17128
rect 17218 17076 17224 17128
rect 17276 17116 17282 17128
rect 18141 17119 18199 17125
rect 18141 17116 18153 17119
rect 17276 17088 18153 17116
rect 17276 17076 17282 17088
rect 18141 17085 18153 17088
rect 18187 17085 18199 17119
rect 18141 17079 18199 17085
rect 7837 17051 7895 17057
rect 7837 17048 7849 17051
rect 5736 17020 7849 17048
rect 5629 17011 5687 17017
rect 7837 17017 7849 17020
rect 7883 17017 7895 17051
rect 7837 17011 7895 17017
rect 11885 17051 11943 17057
rect 11885 17017 11897 17051
rect 11931 17048 11943 17051
rect 12618 17048 12624 17060
rect 11931 17020 12624 17048
rect 11931 17017 11943 17020
rect 11885 17011 11943 17017
rect 12618 17008 12624 17020
rect 12676 17008 12682 17060
rect 15746 17008 15752 17060
rect 15804 17048 15810 17060
rect 18156 17048 18184 17079
rect 18598 17076 18604 17128
rect 18656 17076 18662 17128
rect 19426 17116 19432 17128
rect 19387 17088 19432 17116
rect 19426 17076 19432 17088
rect 19484 17076 19490 17128
rect 19909 17116 19937 17147
rect 20162 17144 20168 17159
rect 20220 17144 20226 17196
rect 20916 17193 20944 17224
rect 21192 17193 21220 17292
rect 22462 17280 22468 17332
rect 22520 17320 22526 17332
rect 22557 17323 22615 17329
rect 22557 17320 22569 17323
rect 22520 17292 22569 17320
rect 22520 17280 22526 17292
rect 22557 17289 22569 17292
rect 22603 17289 22615 17323
rect 26970 17320 26976 17332
rect 26931 17292 26976 17320
rect 22557 17283 22615 17289
rect 26970 17280 26976 17292
rect 27028 17280 27034 17332
rect 28350 17280 28356 17332
rect 28408 17320 28414 17332
rect 29273 17323 29331 17329
rect 29273 17320 29285 17323
rect 28408 17292 29285 17320
rect 28408 17280 28414 17292
rect 29273 17289 29285 17292
rect 29319 17289 29331 17323
rect 29273 17283 29331 17289
rect 31846 17280 31852 17332
rect 31904 17320 31910 17332
rect 31904 17292 33824 17320
rect 31904 17280 31910 17292
rect 24949 17255 25007 17261
rect 24949 17221 24961 17255
rect 24995 17252 25007 17255
rect 28810 17252 28816 17264
rect 24995 17224 27200 17252
rect 24995 17221 25007 17224
rect 24949 17215 25007 17221
rect 20809 17187 20867 17193
rect 20723 17159 20821 17187
rect 20723 17128 20751 17159
rect 20809 17153 20821 17159
rect 20855 17153 20867 17187
rect 20809 17147 20867 17153
rect 20901 17187 20959 17193
rect 20901 17153 20913 17187
rect 20947 17153 20959 17187
rect 20901 17147 20959 17153
rect 20993 17187 21051 17193
rect 20993 17153 21005 17187
rect 21039 17153 21051 17187
rect 20993 17147 21051 17153
rect 21177 17187 21235 17193
rect 21177 17153 21189 17187
rect 21223 17153 21235 17187
rect 21177 17147 21235 17153
rect 19909 17088 20208 17116
rect 20180 17060 20208 17088
rect 20714 17076 20720 17128
rect 20772 17076 20778 17128
rect 19242 17048 19248 17060
rect 15804 17020 17356 17048
rect 18156 17020 19248 17048
rect 15804 17008 15810 17020
rect 4065 16983 4123 16989
rect 4065 16949 4077 16983
rect 4111 16980 4123 16983
rect 5534 16980 5540 16992
rect 4111 16952 5540 16980
rect 4111 16949 4123 16952
rect 4065 16943 4123 16949
rect 5534 16940 5540 16952
rect 5592 16940 5598 16992
rect 8202 16940 8208 16992
rect 8260 16980 8266 16992
rect 8481 16983 8539 16989
rect 8481 16980 8493 16983
rect 8260 16952 8493 16980
rect 8260 16940 8266 16952
rect 8481 16949 8493 16952
rect 8527 16949 8539 16983
rect 14918 16980 14924 16992
rect 14879 16952 14924 16980
rect 8481 16943 8539 16949
rect 14918 16940 14924 16952
rect 14976 16940 14982 16992
rect 16022 16980 16028 16992
rect 15983 16952 16028 16980
rect 16022 16940 16028 16952
rect 16080 16940 16086 16992
rect 17034 16940 17040 16992
rect 17092 16980 17098 16992
rect 17221 16983 17279 16989
rect 17221 16980 17233 16983
rect 17092 16952 17233 16980
rect 17092 16940 17098 16952
rect 17221 16949 17233 16952
rect 17267 16949 17279 16983
rect 17328 16980 17356 17020
rect 19242 17008 19248 17020
rect 19300 17008 19306 17060
rect 20162 17008 20168 17060
rect 20220 17048 20226 17060
rect 21008 17048 21036 17147
rect 21450 17144 21456 17196
rect 21508 17184 21514 17196
rect 21913 17187 21971 17193
rect 21913 17184 21925 17187
rect 21508 17156 21925 17184
rect 21508 17144 21514 17156
rect 21913 17153 21925 17156
rect 21959 17153 21971 17187
rect 23290 17184 23296 17196
rect 23251 17156 23296 17184
rect 21913 17147 21971 17153
rect 23290 17144 23296 17156
rect 23348 17144 23354 17196
rect 23569 17187 23627 17193
rect 23569 17153 23581 17187
rect 23615 17184 23627 17187
rect 24581 17187 24639 17193
rect 24581 17184 24593 17187
rect 23615 17156 24593 17184
rect 23615 17153 23627 17156
rect 23569 17147 23627 17153
rect 24581 17153 24593 17156
rect 24627 17184 24639 17187
rect 24670 17184 24676 17196
rect 24627 17156 24676 17184
rect 24627 17153 24639 17156
rect 24581 17147 24639 17153
rect 24670 17144 24676 17156
rect 24728 17144 24734 17196
rect 24765 17187 24823 17193
rect 24765 17153 24777 17187
rect 24811 17184 24823 17187
rect 25590 17184 25596 17196
rect 24811 17156 25596 17184
rect 24811 17153 24823 17156
rect 24765 17147 24823 17153
rect 25590 17144 25596 17156
rect 25648 17144 25654 17196
rect 25869 17187 25927 17193
rect 25869 17153 25881 17187
rect 25915 17153 25927 17187
rect 26142 17184 26148 17196
rect 26103 17156 26148 17184
rect 25869 17147 25927 17153
rect 21634 17076 21640 17128
rect 21692 17116 21698 17128
rect 22370 17116 22376 17128
rect 21692 17088 22376 17116
rect 21692 17076 21698 17088
rect 22370 17076 22376 17088
rect 22428 17076 22434 17128
rect 25884 17116 25912 17147
rect 26142 17144 26148 17156
rect 26200 17144 26206 17196
rect 27172 17193 27200 17224
rect 27908 17224 28816 17252
rect 27157 17187 27215 17193
rect 27157 17153 27169 17187
rect 27203 17153 27215 17187
rect 27157 17147 27215 17153
rect 26326 17116 26332 17128
rect 25884 17088 26332 17116
rect 26326 17076 26332 17088
rect 26384 17076 26390 17128
rect 27246 17076 27252 17128
rect 27304 17116 27310 17128
rect 27908 17125 27936 17224
rect 28810 17212 28816 17224
rect 28868 17252 28874 17264
rect 30650 17252 30656 17264
rect 28868 17224 30656 17252
rect 28868 17212 28874 17224
rect 28160 17187 28218 17193
rect 28160 17153 28172 17187
rect 28206 17184 28218 17187
rect 28626 17184 28632 17196
rect 28206 17156 28632 17184
rect 28206 17153 28218 17156
rect 28160 17147 28218 17153
rect 28626 17144 28632 17156
rect 28684 17144 28690 17196
rect 29748 17193 29776 17224
rect 30650 17212 30656 17224
rect 30708 17212 30714 17264
rect 32309 17255 32367 17261
rect 32309 17221 32321 17255
rect 32355 17252 32367 17255
rect 33410 17252 33416 17264
rect 32355 17224 33416 17252
rect 32355 17221 32367 17224
rect 32309 17215 32367 17221
rect 33410 17212 33416 17224
rect 33468 17212 33474 17264
rect 29733 17187 29791 17193
rect 29733 17153 29745 17187
rect 29779 17153 29791 17187
rect 29733 17147 29791 17153
rect 29822 17144 29828 17196
rect 29880 17184 29886 17196
rect 29989 17187 30047 17193
rect 29989 17184 30001 17187
rect 29880 17156 30001 17184
rect 29880 17144 29886 17156
rect 29989 17153 30001 17156
rect 30035 17153 30047 17187
rect 29989 17147 30047 17153
rect 31294 17144 31300 17196
rect 31352 17184 31358 17196
rect 33796 17193 33824 17292
rect 34146 17212 34152 17264
rect 34204 17252 34210 17264
rect 34946 17255 35004 17261
rect 34946 17252 34958 17255
rect 34204 17224 34958 17252
rect 34204 17212 34210 17224
rect 34946 17221 34958 17224
rect 34992 17221 35004 17255
rect 34946 17215 35004 17221
rect 32125 17187 32183 17193
rect 32125 17184 32137 17187
rect 31352 17156 32137 17184
rect 31352 17144 31358 17156
rect 32125 17153 32137 17156
rect 32171 17153 32183 17187
rect 32125 17147 32183 17153
rect 33137 17187 33195 17193
rect 33137 17153 33149 17187
rect 33183 17153 33195 17187
rect 33137 17147 33195 17153
rect 33781 17187 33839 17193
rect 33781 17153 33793 17187
rect 33827 17153 33839 17187
rect 33781 17147 33839 17153
rect 27893 17119 27951 17125
rect 27893 17116 27905 17119
rect 27304 17088 27905 17116
rect 27304 17076 27310 17088
rect 27893 17085 27905 17088
rect 27939 17085 27951 17119
rect 27893 17079 27951 17085
rect 31938 17076 31944 17128
rect 31996 17116 32002 17128
rect 33152 17116 33180 17147
rect 31996 17088 33180 17116
rect 31996 17076 32002 17088
rect 34422 17076 34428 17128
rect 34480 17116 34486 17128
rect 34701 17119 34759 17125
rect 34701 17116 34713 17119
rect 34480 17088 34713 17116
rect 34480 17076 34486 17088
rect 34701 17085 34713 17088
rect 34747 17085 34759 17119
rect 34701 17079 34759 17085
rect 20220 17020 21036 17048
rect 20220 17008 20226 17020
rect 25038 17008 25044 17060
rect 25096 17048 25102 17060
rect 26053 17051 26111 17057
rect 26053 17048 26065 17051
rect 25096 17020 26065 17048
rect 25096 17008 25102 17020
rect 26053 17017 26065 17020
rect 26099 17048 26111 17051
rect 26142 17048 26148 17060
rect 26099 17020 26148 17048
rect 26099 17017 26111 17020
rect 26053 17011 26111 17017
rect 26142 17008 26148 17020
rect 26200 17008 26206 17060
rect 32953 17051 33011 17057
rect 32953 17017 32965 17051
rect 32999 17048 33011 17051
rect 33962 17048 33968 17060
rect 32999 17020 33968 17048
rect 32999 17017 33011 17020
rect 32953 17011 33011 17017
rect 33962 17008 33968 17020
rect 34020 17008 34026 17060
rect 20070 16980 20076 16992
rect 17328 16952 20076 16980
rect 17221 16943 17279 16949
rect 20070 16940 20076 16952
rect 20128 16940 20134 16992
rect 20530 16980 20536 16992
rect 20491 16952 20536 16980
rect 20530 16940 20536 16952
rect 20588 16940 20594 16992
rect 25590 16940 25596 16992
rect 25648 16980 25654 16992
rect 25685 16983 25743 16989
rect 25685 16980 25697 16983
rect 25648 16952 25697 16980
rect 25648 16940 25654 16952
rect 25685 16949 25697 16952
rect 25731 16949 25743 16983
rect 25685 16943 25743 16949
rect 30834 16940 30840 16992
rect 30892 16980 30898 16992
rect 31113 16983 31171 16989
rect 31113 16980 31125 16983
rect 30892 16952 31125 16980
rect 30892 16940 30898 16952
rect 31113 16949 31125 16952
rect 31159 16949 31171 16983
rect 32490 16980 32496 16992
rect 32451 16952 32496 16980
rect 31113 16943 31171 16949
rect 32490 16940 32496 16952
rect 32548 16940 32554 16992
rect 33597 16983 33655 16989
rect 33597 16949 33609 16983
rect 33643 16980 33655 16983
rect 33778 16980 33784 16992
rect 33643 16952 33784 16980
rect 33643 16949 33655 16952
rect 33597 16943 33655 16949
rect 33778 16940 33784 16952
rect 33836 16940 33842 16992
rect 34514 16940 34520 16992
rect 34572 16980 34578 16992
rect 36081 16983 36139 16989
rect 36081 16980 36093 16983
rect 34572 16952 36093 16980
rect 34572 16940 34578 16952
rect 36081 16949 36093 16952
rect 36127 16949 36139 16983
rect 36081 16943 36139 16949
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 7374 16776 7380 16788
rect 7335 16748 7380 16776
rect 7374 16736 7380 16748
rect 7432 16736 7438 16788
rect 9030 16776 9036 16788
rect 8312 16748 9036 16776
rect 5169 16711 5227 16717
rect 5169 16677 5181 16711
rect 5215 16677 5227 16711
rect 8312 16708 8340 16748
rect 9030 16736 9036 16748
rect 9088 16736 9094 16788
rect 9306 16776 9312 16788
rect 9267 16748 9312 16776
rect 9306 16736 9312 16748
rect 9364 16736 9370 16788
rect 13722 16776 13728 16788
rect 11256 16748 13728 16776
rect 8846 16708 8852 16720
rect 5169 16671 5227 16677
rect 6564 16680 8340 16708
rect 8404 16680 8852 16708
rect 2866 16600 2872 16652
rect 2924 16640 2930 16652
rect 3786 16640 3792 16652
rect 2924 16612 3792 16640
rect 2924 16600 2930 16612
rect 3786 16600 3792 16612
rect 3844 16600 3850 16652
rect 1854 16572 1860 16584
rect 1767 16544 1860 16572
rect 1854 16532 1860 16544
rect 1912 16572 1918 16584
rect 2682 16572 2688 16584
rect 1912 16544 2688 16572
rect 1912 16532 1918 16544
rect 2682 16532 2688 16544
rect 2740 16532 2746 16584
rect 4062 16581 4068 16584
rect 4056 16572 4068 16581
rect 4023 16544 4068 16572
rect 4056 16535 4068 16544
rect 4062 16532 4068 16535
rect 4120 16532 4126 16584
rect 5184 16572 5212 16671
rect 6564 16649 6592 16680
rect 6549 16643 6607 16649
rect 6549 16609 6561 16643
rect 6595 16609 6607 16643
rect 6549 16603 6607 16609
rect 8404 16581 8432 16680
rect 8846 16668 8852 16680
rect 8904 16668 8910 16720
rect 10686 16668 10692 16720
rect 10744 16708 10750 16720
rect 11256 16708 11284 16748
rect 13722 16736 13728 16748
rect 13780 16736 13786 16788
rect 15010 16736 15016 16788
rect 15068 16736 15074 16788
rect 24765 16779 24823 16785
rect 19260 16748 22094 16776
rect 14734 16708 14740 16720
rect 10744 16680 11284 16708
rect 10744 16668 10750 16680
rect 11256 16640 11284 16680
rect 13004 16680 14740 16708
rect 11164 16612 11284 16640
rect 7193 16575 7251 16581
rect 7193 16572 7205 16575
rect 5184 16544 7205 16572
rect 7193 16541 7205 16544
rect 7239 16541 7251 16575
rect 7193 16535 7251 16541
rect 8205 16575 8263 16581
rect 8205 16541 8217 16575
rect 8251 16541 8263 16575
rect 8205 16535 8263 16541
rect 8389 16575 8447 16581
rect 8389 16541 8401 16575
rect 8435 16541 8447 16575
rect 8389 16535 8447 16541
rect 2124 16507 2182 16513
rect 2124 16473 2136 16507
rect 2170 16504 2182 16507
rect 5718 16504 5724 16516
rect 2170 16476 5724 16504
rect 2170 16473 2182 16476
rect 2124 16467 2182 16473
rect 5718 16464 5724 16476
rect 5776 16464 5782 16516
rect 5994 16464 6000 16516
rect 6052 16504 6058 16516
rect 6181 16507 6239 16513
rect 6181 16504 6193 16507
rect 6052 16476 6193 16504
rect 6052 16464 6058 16476
rect 6181 16473 6193 16476
rect 6227 16473 6239 16507
rect 6181 16467 6239 16473
rect 6365 16507 6423 16513
rect 6365 16473 6377 16507
rect 6411 16473 6423 16507
rect 7006 16504 7012 16516
rect 6967 16476 7012 16504
rect 6365 16467 6423 16473
rect 3237 16439 3295 16445
rect 3237 16405 3249 16439
rect 3283 16436 3295 16439
rect 5074 16436 5080 16448
rect 3283 16408 5080 16436
rect 3283 16405 3295 16408
rect 3237 16399 3295 16405
rect 5074 16396 5080 16408
rect 5132 16396 5138 16448
rect 5626 16396 5632 16448
rect 5684 16436 5690 16448
rect 6380 16436 6408 16467
rect 7006 16464 7012 16476
rect 7064 16464 7070 16516
rect 5684 16408 6408 16436
rect 7024 16436 7052 16464
rect 7190 16436 7196 16448
rect 7024 16408 7196 16436
rect 5684 16396 5690 16408
rect 7190 16396 7196 16408
rect 7248 16396 7254 16448
rect 8220 16436 8248 16535
rect 10962 16532 10968 16584
rect 11020 16581 11026 16584
rect 11164 16581 11192 16612
rect 11330 16600 11336 16652
rect 11388 16640 11394 16652
rect 11388 16612 11468 16640
rect 11388 16600 11394 16612
rect 11020 16575 11069 16581
rect 11020 16541 11023 16575
rect 11057 16541 11069 16575
rect 11020 16535 11069 16541
rect 11146 16575 11204 16581
rect 11146 16541 11158 16575
rect 11192 16541 11204 16575
rect 11146 16535 11204 16541
rect 11020 16532 11026 16535
rect 11238 16532 11244 16584
rect 11296 16581 11302 16584
rect 11440 16581 11468 16612
rect 11296 16572 11304 16581
rect 11425 16575 11483 16581
rect 11296 16544 11341 16572
rect 11296 16535 11304 16544
rect 11425 16541 11437 16575
rect 11471 16541 11483 16575
rect 11425 16535 11483 16541
rect 11296 16532 11302 16535
rect 8297 16507 8355 16513
rect 8297 16473 8309 16507
rect 8343 16504 8355 16507
rect 8938 16504 8944 16516
rect 8343 16476 8944 16504
rect 8343 16473 8355 16476
rect 8297 16467 8355 16473
rect 8938 16464 8944 16476
rect 8996 16464 9002 16516
rect 9122 16504 9128 16516
rect 9083 16476 9128 16504
rect 9122 16464 9128 16476
rect 9180 16464 9186 16516
rect 10980 16504 11008 16532
rect 13004 16504 13032 16680
rect 14734 16668 14740 16680
rect 14792 16708 14798 16720
rect 14792 16680 14872 16708
rect 14792 16668 14798 16680
rect 14844 16640 14872 16680
rect 14844 16612 14964 16640
rect 13078 16532 13084 16584
rect 13136 16550 13142 16584
rect 13173 16575 13231 16581
rect 13173 16550 13185 16575
rect 13136 16541 13185 16550
rect 13219 16541 13231 16575
rect 13136 16535 13231 16541
rect 13262 16572 13320 16578
rect 13262 16562 13274 16572
rect 13308 16562 13320 16572
rect 13357 16575 13415 16581
rect 13136 16532 13216 16535
rect 13096 16522 13216 16532
rect 13262 16510 13268 16562
rect 13320 16510 13326 16562
rect 13357 16541 13369 16575
rect 13403 16541 13415 16575
rect 13357 16535 13415 16541
rect 13553 16575 13611 16581
rect 13553 16541 13565 16575
rect 13599 16572 13611 16575
rect 13998 16572 14004 16584
rect 13599 16544 14004 16572
rect 13599 16541 13611 16544
rect 13553 16535 13611 16541
rect 10980 16476 13032 16504
rect 9398 16436 9404 16448
rect 8220 16408 9404 16436
rect 9398 16396 9404 16408
rect 9456 16396 9462 16448
rect 10781 16439 10839 16445
rect 10781 16405 10793 16439
rect 10827 16436 10839 16439
rect 10962 16436 10968 16448
rect 10827 16408 10968 16436
rect 10827 16405 10839 16408
rect 10781 16399 10839 16405
rect 10962 16396 10968 16408
rect 11020 16396 11026 16448
rect 12897 16439 12955 16445
rect 12897 16405 12909 16439
rect 12943 16436 12955 16439
rect 13078 16436 13084 16448
rect 12943 16408 13084 16436
rect 12943 16405 12955 16408
rect 12897 16399 12955 16405
rect 13078 16396 13084 16408
rect 13136 16396 13142 16448
rect 13170 16396 13176 16448
rect 13228 16436 13234 16448
rect 13372 16436 13400 16535
rect 13998 16532 14004 16544
rect 14056 16572 14062 16584
rect 14936 16581 14964 16612
rect 15028 16581 15056 16736
rect 15562 16668 15568 16720
rect 15620 16708 15626 16720
rect 15620 16680 18000 16708
rect 15620 16668 15626 16680
rect 17126 16640 17132 16652
rect 15856 16612 17132 16640
rect 14921 16575 14979 16581
rect 14056 16544 14872 16572
rect 14056 16532 14062 16544
rect 14844 16504 14872 16544
rect 14921 16541 14933 16575
rect 14967 16541 14979 16575
rect 14921 16535 14979 16541
rect 15013 16575 15071 16581
rect 15013 16541 15025 16575
rect 15059 16541 15071 16575
rect 15013 16535 15071 16541
rect 15102 16532 15108 16584
rect 15160 16572 15166 16584
rect 15160 16544 15205 16572
rect 15160 16532 15166 16544
rect 15286 16532 15292 16584
rect 15344 16572 15350 16584
rect 15746 16572 15752 16584
rect 15344 16544 15389 16572
rect 15707 16544 15752 16572
rect 15344 16532 15350 16544
rect 15746 16532 15752 16544
rect 15804 16532 15810 16584
rect 15856 16504 15884 16612
rect 17126 16600 17132 16612
rect 17184 16640 17190 16652
rect 17184 16612 17264 16640
rect 17184 16600 17190 16612
rect 16850 16572 16856 16584
rect 16811 16544 16856 16572
rect 16850 16532 16856 16544
rect 16908 16532 16914 16584
rect 16945 16575 17003 16581
rect 16945 16541 16957 16575
rect 16991 16541 17003 16575
rect 16945 16535 17003 16541
rect 14844 16476 15884 16504
rect 16960 16504 16988 16535
rect 17034 16532 17040 16584
rect 17092 16581 17098 16584
rect 17236 16581 17264 16612
rect 17092 16572 17100 16581
rect 17221 16575 17279 16581
rect 17092 16544 17137 16572
rect 17092 16535 17100 16544
rect 17221 16541 17233 16575
rect 17267 16541 17279 16575
rect 17221 16535 17279 16541
rect 17092 16532 17098 16535
rect 17586 16532 17592 16584
rect 17644 16572 17650 16584
rect 17972 16581 18000 16680
rect 18138 16668 18144 16720
rect 18196 16708 18202 16720
rect 18196 16680 18276 16708
rect 18196 16668 18202 16680
rect 17865 16575 17923 16581
rect 17865 16572 17877 16575
rect 17644 16544 17877 16572
rect 17644 16532 17650 16544
rect 17865 16541 17877 16544
rect 17911 16541 17923 16575
rect 17865 16535 17923 16541
rect 17957 16575 18015 16581
rect 17957 16541 17969 16575
rect 18003 16541 18015 16575
rect 18138 16572 18144 16584
rect 18099 16544 18144 16572
rect 17957 16535 18015 16541
rect 18138 16532 18144 16544
rect 18196 16532 18202 16584
rect 18248 16581 18276 16680
rect 19260 16649 19288 16748
rect 21450 16708 21456 16720
rect 21411 16680 21456 16708
rect 21450 16668 21456 16680
rect 21508 16668 21514 16720
rect 19245 16643 19303 16649
rect 19245 16609 19257 16643
rect 19291 16609 19303 16643
rect 22066 16640 22094 16748
rect 24765 16745 24777 16779
rect 24811 16776 24823 16779
rect 25038 16776 25044 16788
rect 24811 16748 25044 16776
rect 24811 16745 24823 16748
rect 24765 16739 24823 16745
rect 25038 16736 25044 16748
rect 25096 16736 25102 16788
rect 29733 16779 29791 16785
rect 29733 16745 29745 16779
rect 29779 16776 29791 16779
rect 29822 16776 29828 16788
rect 29779 16748 29828 16776
rect 29779 16745 29791 16748
rect 29733 16739 29791 16745
rect 29822 16736 29828 16748
rect 29880 16736 29886 16788
rect 32490 16736 32496 16788
rect 32548 16776 32554 16788
rect 35802 16776 35808 16788
rect 32548 16748 35808 16776
rect 32548 16736 32554 16748
rect 35802 16736 35808 16748
rect 35860 16736 35866 16788
rect 31662 16708 31668 16720
rect 24412 16680 24992 16708
rect 31623 16680 31668 16708
rect 22186 16640 22192 16652
rect 19245 16603 19303 16609
rect 21284 16612 21772 16640
rect 22066 16612 22192 16640
rect 18233 16575 18291 16581
rect 18233 16541 18245 16575
rect 18279 16541 18291 16575
rect 18233 16535 18291 16541
rect 19512 16575 19570 16581
rect 19512 16541 19524 16575
rect 19558 16572 19570 16575
rect 20530 16572 20536 16584
rect 19558 16544 20536 16572
rect 19558 16541 19570 16544
rect 19512 16535 19570 16541
rect 20530 16532 20536 16544
rect 20588 16532 20594 16584
rect 20622 16532 20628 16584
rect 20680 16572 20686 16584
rect 20806 16572 20812 16584
rect 20680 16544 20812 16572
rect 20680 16532 20686 16544
rect 20806 16532 20812 16544
rect 20864 16532 20870 16584
rect 17604 16504 17632 16532
rect 21284 16504 21312 16612
rect 21744 16584 21772 16612
rect 22186 16600 22192 16612
rect 22244 16640 22250 16652
rect 22465 16643 22523 16649
rect 22465 16640 22477 16643
rect 22244 16612 22477 16640
rect 22244 16600 22250 16612
rect 22465 16609 22477 16612
rect 22511 16609 22523 16643
rect 22465 16603 22523 16609
rect 21634 16572 21640 16584
rect 21595 16544 21640 16572
rect 21634 16532 21640 16544
rect 21692 16532 21698 16584
rect 21726 16532 21732 16584
rect 21784 16572 21790 16584
rect 21913 16575 21971 16581
rect 21784 16544 21877 16572
rect 21784 16532 21790 16544
rect 21913 16541 21925 16575
rect 21959 16541 21971 16575
rect 21913 16535 21971 16541
rect 22005 16575 22063 16581
rect 22005 16541 22017 16575
rect 22051 16572 22063 16575
rect 23474 16572 23480 16584
rect 22051 16544 23480 16572
rect 22051 16541 22063 16544
rect 22005 16535 22063 16541
rect 16960 16476 17632 16504
rect 17972 16476 21312 16504
rect 21928 16504 21956 16535
rect 23474 16532 23480 16544
rect 23532 16532 23538 16584
rect 24412 16572 24440 16680
rect 24857 16643 24915 16649
rect 24857 16609 24869 16643
rect 24903 16609 24915 16643
rect 24857 16603 24915 16609
rect 24578 16572 24584 16584
rect 23584 16544 24440 16572
rect 24539 16544 24584 16572
rect 22554 16504 22560 16516
rect 21928 16476 22560 16504
rect 17972 16448 18000 16476
rect 22554 16464 22560 16476
rect 22612 16464 22618 16516
rect 22732 16507 22790 16513
rect 22732 16473 22744 16507
rect 22778 16504 22790 16507
rect 23290 16504 23296 16516
rect 22778 16476 23296 16504
rect 22778 16473 22790 16476
rect 22732 16467 22790 16473
rect 23290 16464 23296 16476
rect 23348 16464 23354 16516
rect 23382 16464 23388 16516
rect 23440 16504 23446 16516
rect 23584 16504 23612 16544
rect 24578 16532 24584 16544
rect 24636 16532 24642 16584
rect 24872 16504 24900 16603
rect 24964 16572 24992 16680
rect 31662 16668 31668 16680
rect 31720 16668 31726 16720
rect 33781 16711 33839 16717
rect 33781 16677 33793 16711
rect 33827 16708 33839 16711
rect 33827 16680 33916 16708
rect 33827 16677 33839 16680
rect 33781 16671 33839 16677
rect 26053 16643 26111 16649
rect 26053 16609 26065 16643
rect 26099 16640 26111 16643
rect 27062 16640 27068 16652
rect 26099 16612 27068 16640
rect 26099 16609 26111 16612
rect 26053 16603 26111 16609
rect 27062 16600 27068 16612
rect 27120 16600 27126 16652
rect 27246 16640 27252 16652
rect 27207 16612 27252 16640
rect 27246 16600 27252 16612
rect 27304 16600 27310 16652
rect 30377 16643 30435 16649
rect 30377 16609 30389 16643
rect 30423 16640 30435 16643
rect 30466 16640 30472 16652
rect 30423 16612 30472 16640
rect 30423 16609 30435 16612
rect 30377 16603 30435 16609
rect 30466 16600 30472 16612
rect 30524 16600 30530 16652
rect 30834 16640 30840 16652
rect 30795 16612 30840 16640
rect 30834 16600 30840 16612
rect 30892 16600 30898 16652
rect 32493 16643 32551 16649
rect 32493 16609 32505 16643
rect 32539 16640 32551 16643
rect 33321 16643 33379 16649
rect 32539 16612 33272 16640
rect 32539 16609 32551 16612
rect 32493 16603 32551 16609
rect 25869 16575 25927 16581
rect 25869 16572 25881 16575
rect 24964 16544 25881 16572
rect 25869 16541 25881 16544
rect 25915 16541 25927 16575
rect 25869 16535 25927 16541
rect 26142 16532 26148 16584
rect 26200 16572 26206 16584
rect 29914 16572 29920 16584
rect 26200 16544 29776 16572
rect 29875 16544 29920 16572
rect 26200 16532 26206 16544
rect 23440 16476 23612 16504
rect 23860 16476 24900 16504
rect 27516 16507 27574 16513
rect 23440 16464 23446 16476
rect 13228 16408 13400 16436
rect 13228 16396 13234 16408
rect 13446 16396 13452 16448
rect 13504 16436 13510 16448
rect 14645 16439 14703 16445
rect 14645 16436 14657 16439
rect 13504 16408 14657 16436
rect 13504 16396 13510 16408
rect 14645 16405 14657 16408
rect 14691 16405 14703 16439
rect 14645 16399 14703 16405
rect 15470 16396 15476 16448
rect 15528 16436 15534 16448
rect 15933 16439 15991 16445
rect 15933 16436 15945 16439
rect 15528 16408 15945 16436
rect 15528 16396 15534 16408
rect 15933 16405 15945 16408
rect 15979 16436 15991 16439
rect 16206 16436 16212 16448
rect 15979 16408 16212 16436
rect 15979 16405 15991 16408
rect 15933 16399 15991 16405
rect 16206 16396 16212 16408
rect 16264 16396 16270 16448
rect 16390 16396 16396 16448
rect 16448 16436 16454 16448
rect 16577 16439 16635 16445
rect 16577 16436 16589 16439
rect 16448 16408 16589 16436
rect 16448 16396 16454 16408
rect 16577 16405 16589 16408
rect 16623 16405 16635 16439
rect 16577 16399 16635 16405
rect 17034 16396 17040 16448
rect 17092 16436 17098 16448
rect 17681 16439 17739 16445
rect 17681 16436 17693 16439
rect 17092 16408 17693 16436
rect 17092 16396 17098 16408
rect 17681 16405 17693 16408
rect 17727 16405 17739 16439
rect 17681 16399 17739 16405
rect 17954 16396 17960 16448
rect 18012 16396 18018 16448
rect 20070 16396 20076 16448
rect 20128 16436 20134 16448
rect 20625 16439 20683 16445
rect 20625 16436 20637 16439
rect 20128 16408 20637 16436
rect 20128 16396 20134 16408
rect 20625 16405 20637 16408
rect 20671 16405 20683 16439
rect 20625 16399 20683 16405
rect 23106 16396 23112 16448
rect 23164 16436 23170 16448
rect 23400 16436 23428 16464
rect 23860 16445 23888 16476
rect 27516 16473 27528 16507
rect 27562 16504 27574 16507
rect 27614 16504 27620 16516
rect 27562 16476 27620 16504
rect 27562 16473 27574 16476
rect 27516 16467 27574 16473
rect 27614 16464 27620 16476
rect 27672 16464 27678 16516
rect 23164 16408 23428 16436
rect 23845 16439 23903 16445
rect 23164 16396 23170 16408
rect 23845 16405 23857 16439
rect 23891 16405 23903 16439
rect 24394 16436 24400 16448
rect 24355 16408 24400 16436
rect 23845 16399 23903 16405
rect 24394 16396 24400 16408
rect 24452 16396 24458 16448
rect 28350 16396 28356 16448
rect 28408 16436 28414 16448
rect 28629 16439 28687 16445
rect 28629 16436 28641 16439
rect 28408 16408 28641 16436
rect 28408 16396 28414 16408
rect 28629 16405 28641 16408
rect 28675 16405 28687 16439
rect 29748 16436 29776 16544
rect 29914 16532 29920 16544
rect 29972 16532 29978 16584
rect 30561 16575 30619 16581
rect 30561 16541 30573 16575
rect 30607 16541 30619 16575
rect 30742 16572 30748 16584
rect 30703 16544 30748 16572
rect 30561 16535 30619 16541
rect 30576 16504 30604 16535
rect 30742 16532 30748 16544
rect 30800 16532 30806 16584
rect 30926 16532 30932 16584
rect 30984 16572 30990 16584
rect 31294 16572 31300 16584
rect 30984 16544 31300 16572
rect 30984 16532 30990 16544
rect 31294 16532 31300 16544
rect 31352 16572 31358 16584
rect 32309 16575 32367 16581
rect 31352 16544 31708 16572
rect 31352 16532 31358 16544
rect 31680 16516 31708 16544
rect 32309 16541 32321 16575
rect 32355 16572 32367 16575
rect 33042 16572 33048 16584
rect 32355 16544 33048 16572
rect 32355 16541 32367 16544
rect 32309 16535 32367 16541
rect 33042 16532 33048 16544
rect 33100 16532 33106 16584
rect 33244 16572 33272 16612
rect 33321 16609 33333 16643
rect 33367 16640 33379 16643
rect 33594 16640 33600 16652
rect 33367 16612 33600 16640
rect 33367 16609 33379 16612
rect 33321 16603 33379 16609
rect 33594 16600 33600 16612
rect 33652 16600 33658 16652
rect 33888 16640 33916 16680
rect 34790 16640 34796 16652
rect 33888 16612 34796 16640
rect 34790 16600 34796 16612
rect 34848 16600 34854 16652
rect 33965 16575 34023 16581
rect 33965 16572 33977 16575
rect 33244 16548 33640 16572
rect 33888 16548 33977 16572
rect 33244 16544 33977 16548
rect 33612 16520 33916 16544
rect 33965 16541 33977 16544
rect 34011 16541 34023 16575
rect 33965 16535 34023 16541
rect 31110 16504 31116 16516
rect 30576 16476 31116 16504
rect 31110 16464 31116 16476
rect 31168 16464 31174 16516
rect 31478 16504 31484 16516
rect 31439 16476 31484 16504
rect 31478 16464 31484 16476
rect 31536 16464 31542 16516
rect 31662 16464 31668 16516
rect 31720 16464 31726 16516
rect 32122 16504 32128 16516
rect 32083 16476 32128 16504
rect 32122 16464 32128 16476
rect 32180 16464 32186 16516
rect 32398 16464 32404 16516
rect 32456 16504 32462 16516
rect 32953 16507 33011 16513
rect 32953 16504 32965 16507
rect 32456 16476 32965 16504
rect 32456 16464 32462 16476
rect 32953 16473 32965 16476
rect 32999 16473 33011 16507
rect 32953 16467 33011 16473
rect 33137 16507 33195 16513
rect 33137 16473 33149 16507
rect 33183 16473 33195 16507
rect 33137 16467 33195 16473
rect 30742 16436 30748 16448
rect 29748 16408 30748 16436
rect 28629 16399 28687 16405
rect 30742 16396 30748 16408
rect 30800 16396 30806 16448
rect 31754 16396 31760 16448
rect 31812 16436 31818 16448
rect 32858 16436 32864 16448
rect 31812 16408 32864 16436
rect 31812 16396 31818 16408
rect 32858 16396 32864 16408
rect 32916 16396 32922 16448
rect 33152 16436 33180 16467
rect 34698 16464 34704 16516
rect 34756 16504 34762 16516
rect 35069 16507 35127 16513
rect 35069 16504 35081 16507
rect 34756 16476 35081 16504
rect 34756 16464 34762 16476
rect 35069 16473 35081 16476
rect 35115 16473 35127 16507
rect 35069 16467 35127 16473
rect 33686 16436 33692 16448
rect 33152 16408 33692 16436
rect 33686 16396 33692 16408
rect 33744 16396 33750 16448
rect 34422 16396 34428 16448
rect 34480 16436 34486 16448
rect 36357 16439 36415 16445
rect 36357 16436 36369 16439
rect 34480 16408 36369 16436
rect 34480 16396 34486 16408
rect 36357 16405 36369 16408
rect 36403 16436 36415 16439
rect 36538 16436 36544 16448
rect 36403 16408 36544 16436
rect 36403 16405 36415 16408
rect 36357 16399 36415 16405
rect 36538 16396 36544 16408
rect 36596 16396 36602 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 4065 16235 4123 16241
rect 4065 16201 4077 16235
rect 4111 16232 4123 16235
rect 6733 16235 6791 16241
rect 4111 16204 6592 16232
rect 4111 16201 4123 16204
rect 4065 16195 4123 16201
rect 4706 16124 4712 16176
rect 4764 16164 4770 16176
rect 5629 16167 5687 16173
rect 5629 16164 5641 16167
rect 4764 16136 5641 16164
rect 4764 16124 4770 16136
rect 5629 16133 5641 16136
rect 5675 16133 5687 16167
rect 5810 16164 5816 16176
rect 5771 16136 5816 16164
rect 5629 16127 5687 16133
rect 5810 16124 5816 16136
rect 5868 16124 5874 16176
rect 6564 16173 6592 16204
rect 6733 16201 6745 16235
rect 6779 16232 6791 16235
rect 7834 16232 7840 16244
rect 6779 16204 7840 16232
rect 6779 16201 6791 16204
rect 6733 16195 6791 16201
rect 7834 16192 7840 16204
rect 7892 16192 7898 16244
rect 9122 16192 9128 16244
rect 9180 16232 9186 16244
rect 9309 16235 9367 16241
rect 9309 16232 9321 16235
rect 9180 16204 9321 16232
rect 9180 16192 9186 16204
rect 9309 16201 9321 16204
rect 9355 16201 9367 16235
rect 9309 16195 9367 16201
rect 9398 16192 9404 16244
rect 9456 16232 9462 16244
rect 11790 16232 11796 16244
rect 9456 16204 11796 16232
rect 9456 16192 9462 16204
rect 11790 16192 11796 16204
rect 11848 16192 11854 16244
rect 15657 16235 15715 16241
rect 15657 16201 15669 16235
rect 15703 16232 15715 16235
rect 15930 16232 15936 16244
rect 15703 16204 15936 16232
rect 15703 16201 15715 16204
rect 15657 16195 15715 16201
rect 15930 16192 15936 16204
rect 15988 16192 15994 16244
rect 19981 16235 20039 16241
rect 19981 16201 19993 16235
rect 20027 16232 20039 16235
rect 20162 16232 20168 16244
rect 20027 16204 20168 16232
rect 20027 16201 20039 16204
rect 19981 16195 20039 16201
rect 20162 16192 20168 16204
rect 20220 16192 20226 16244
rect 21726 16192 21732 16244
rect 21784 16232 21790 16244
rect 22002 16232 22008 16244
rect 21784 16204 22008 16232
rect 21784 16192 21790 16204
rect 22002 16192 22008 16204
rect 22060 16192 22066 16244
rect 23474 16232 23480 16244
rect 23216 16204 23480 16232
rect 6549 16167 6607 16173
rect 6549 16133 6561 16167
rect 6595 16133 6607 16167
rect 8018 16164 8024 16176
rect 6549 16127 6607 16133
rect 6748 16136 8024 16164
rect 2682 16096 2688 16108
rect 2643 16068 2688 16096
rect 2682 16056 2688 16068
rect 2740 16056 2746 16108
rect 2952 16099 3010 16105
rect 2952 16065 2964 16099
rect 2998 16096 3010 16099
rect 4985 16099 5043 16105
rect 2998 16068 4936 16096
rect 2998 16065 3010 16068
rect 2952 16059 3010 16065
rect 4798 15892 4804 15904
rect 4759 15864 4804 15892
rect 4798 15852 4804 15864
rect 4856 15852 4862 15904
rect 4908 15892 4936 16068
rect 4985 16065 4997 16099
rect 5031 16065 5043 16099
rect 4985 16059 5043 16065
rect 5000 16028 5028 16059
rect 5350 16056 5356 16108
rect 5408 16096 5414 16108
rect 5445 16099 5503 16105
rect 5445 16096 5457 16099
rect 5408 16068 5457 16096
rect 5408 16056 5414 16068
rect 5445 16065 5457 16068
rect 5491 16096 5503 16099
rect 5994 16096 6000 16108
rect 5491 16068 6000 16096
rect 5491 16065 5503 16068
rect 5445 16059 5503 16065
rect 5994 16056 6000 16068
rect 6052 16056 6058 16108
rect 6362 16096 6368 16108
rect 6323 16068 6368 16096
rect 6362 16056 6368 16068
rect 6420 16056 6426 16108
rect 6270 16028 6276 16040
rect 5000 16000 6276 16028
rect 6270 15988 6276 16000
rect 6328 15988 6334 16040
rect 5074 15920 5080 15972
rect 5132 15960 5138 15972
rect 6638 15960 6644 15972
rect 5132 15932 6644 15960
rect 5132 15920 5138 15932
rect 6638 15920 6644 15932
rect 6696 15920 6702 15972
rect 6748 15892 6776 16136
rect 8018 16124 8024 16136
rect 8076 16124 8082 16176
rect 8202 16173 8208 16176
rect 8196 16164 8208 16173
rect 8163 16136 8208 16164
rect 8196 16127 8208 16136
rect 8202 16124 8208 16127
rect 8260 16124 8266 16176
rect 12618 16164 12624 16176
rect 11072 16136 12624 16164
rect 7374 16096 7380 16108
rect 7335 16068 7380 16096
rect 7374 16056 7380 16068
rect 7432 16056 7438 16108
rect 10597 16099 10655 16105
rect 10597 16065 10609 16099
rect 10643 16065 10655 16099
rect 10597 16059 10655 16065
rect 10686 16099 10744 16105
rect 10686 16065 10698 16099
rect 10732 16065 10744 16099
rect 10686 16059 10744 16065
rect 6822 15988 6828 16040
rect 6880 16028 6886 16040
rect 7929 16031 7987 16037
rect 7929 16028 7941 16031
rect 6880 16000 7941 16028
rect 6880 15988 6886 16000
rect 7929 15997 7941 16000
rect 7975 15997 7987 16031
rect 7929 15991 7987 15997
rect 10502 15988 10508 16040
rect 10560 16028 10566 16040
rect 10612 16028 10640 16059
rect 10560 16000 10640 16028
rect 10560 15988 10566 16000
rect 10704 15972 10732 16059
rect 10778 16056 10784 16108
rect 10836 16105 10842 16108
rect 10836 16096 10844 16105
rect 10965 16099 11023 16105
rect 11072 16099 11100 16136
rect 12618 16124 12624 16136
rect 12676 16124 12682 16176
rect 14544 16167 14602 16173
rect 14544 16133 14556 16167
rect 14590 16164 14602 16167
rect 14918 16164 14924 16176
rect 14590 16136 14924 16164
rect 14590 16133 14602 16136
rect 14544 16127 14602 16133
rect 14918 16124 14924 16136
rect 14976 16124 14982 16176
rect 17310 16164 17316 16176
rect 16776 16136 17316 16164
rect 10836 16068 10881 16096
rect 10836 16059 10844 16068
rect 10965 16065 10977 16099
rect 11011 16071 11100 16099
rect 12428 16099 12486 16105
rect 11011 16065 11023 16071
rect 10965 16059 11023 16065
rect 12428 16065 12440 16099
rect 12474 16096 12486 16099
rect 12710 16096 12716 16108
rect 12474 16068 12716 16096
rect 12474 16065 12486 16068
rect 12428 16059 12486 16065
rect 10836 16056 10842 16059
rect 12710 16056 12716 16068
rect 12768 16056 12774 16108
rect 16776 16105 16804 16136
rect 17310 16124 17316 16136
rect 17368 16124 17374 16176
rect 17862 16124 17868 16176
rect 17920 16164 17926 16176
rect 18693 16167 18751 16173
rect 18693 16164 18705 16167
rect 17920 16136 18705 16164
rect 17920 16124 17926 16136
rect 18693 16133 18705 16136
rect 18739 16133 18751 16167
rect 18693 16127 18751 16133
rect 19334 16124 19340 16176
rect 19392 16164 19398 16176
rect 19613 16167 19671 16173
rect 19613 16164 19625 16167
rect 19392 16136 19625 16164
rect 19392 16124 19398 16136
rect 19613 16133 19625 16136
rect 19659 16133 19671 16167
rect 19613 16127 19671 16133
rect 19797 16167 19855 16173
rect 19797 16133 19809 16167
rect 19843 16164 19855 16167
rect 20070 16164 20076 16176
rect 19843 16136 20076 16164
rect 19843 16133 19855 16136
rect 19797 16127 19855 16133
rect 17034 16105 17040 16108
rect 16761 16099 16819 16105
rect 16761 16065 16773 16099
rect 16807 16065 16819 16099
rect 17028 16096 17040 16105
rect 16995 16068 17040 16096
rect 16761 16059 16819 16065
rect 17028 16059 17040 16068
rect 17034 16056 17040 16059
rect 17092 16056 17098 16108
rect 18601 16099 18659 16105
rect 18601 16096 18613 16099
rect 18156 16068 18613 16096
rect 11146 15988 11152 16040
rect 11204 16028 11210 16040
rect 12161 16031 12219 16037
rect 12161 16028 12173 16031
rect 11204 16000 12173 16028
rect 11204 15988 11210 16000
rect 12161 15997 12173 16000
rect 12207 15997 12219 16031
rect 12161 15991 12219 15997
rect 14277 16031 14335 16037
rect 14277 15997 14289 16031
rect 14323 15997 14335 16031
rect 14277 15991 14335 15997
rect 8864 15932 10456 15960
rect 4908 15864 6776 15892
rect 6914 15852 6920 15904
rect 6972 15892 6978 15904
rect 7193 15895 7251 15901
rect 7193 15892 7205 15895
rect 6972 15864 7205 15892
rect 6972 15852 6978 15864
rect 7193 15861 7205 15864
rect 7239 15861 7251 15895
rect 7193 15855 7251 15861
rect 7282 15852 7288 15904
rect 7340 15892 7346 15904
rect 8864 15892 8892 15932
rect 10318 15892 10324 15904
rect 7340 15864 8892 15892
rect 10279 15864 10324 15892
rect 7340 15852 7346 15864
rect 10318 15852 10324 15864
rect 10376 15852 10382 15904
rect 10428 15892 10456 15932
rect 10686 15920 10692 15972
rect 10744 15920 10750 15972
rect 13446 15960 13452 15972
rect 13372 15932 13452 15960
rect 13372 15892 13400 15932
rect 13446 15920 13452 15932
rect 13504 15920 13510 15972
rect 13538 15892 13544 15904
rect 10428 15864 13400 15892
rect 13499 15864 13544 15892
rect 13538 15852 13544 15864
rect 13596 15852 13602 15904
rect 14292 15892 14320 15991
rect 18156 15969 18184 16068
rect 18601 16065 18613 16068
rect 18647 16065 18659 16099
rect 19628 16096 19656 16127
rect 20070 16124 20076 16136
rect 20128 16124 20134 16176
rect 21913 16167 21971 16173
rect 21913 16164 21925 16167
rect 20548 16136 21925 16164
rect 20548 16096 20576 16136
rect 21913 16133 21925 16136
rect 21959 16164 21971 16167
rect 23106 16164 23112 16176
rect 21959 16136 23112 16164
rect 21959 16133 21971 16136
rect 21913 16127 21971 16133
rect 23106 16124 23112 16136
rect 23164 16124 23170 16176
rect 23216 16173 23244 16204
rect 23474 16192 23480 16204
rect 23532 16232 23538 16244
rect 24670 16232 24676 16244
rect 23532 16204 24676 16232
rect 23532 16192 23538 16204
rect 24670 16192 24676 16204
rect 24728 16192 24734 16244
rect 28626 16192 28632 16244
rect 28684 16232 28690 16244
rect 28813 16235 28871 16241
rect 28813 16232 28825 16235
rect 28684 16204 28825 16232
rect 28684 16192 28690 16204
rect 28813 16201 28825 16204
rect 28859 16201 28871 16235
rect 28813 16195 28871 16201
rect 31478 16192 31484 16244
rect 31536 16232 31542 16244
rect 34057 16235 34115 16241
rect 34057 16232 34069 16235
rect 31536 16204 34069 16232
rect 31536 16192 31542 16204
rect 34057 16201 34069 16204
rect 34103 16201 34115 16235
rect 36357 16235 36415 16241
rect 36357 16232 36369 16235
rect 34057 16195 34115 16201
rect 34532 16204 36369 16232
rect 23201 16167 23259 16173
rect 23201 16133 23213 16167
rect 23247 16133 23259 16167
rect 23201 16127 23259 16133
rect 23385 16167 23443 16173
rect 23385 16133 23397 16167
rect 23431 16164 23443 16167
rect 23842 16164 23848 16176
rect 23431 16136 23848 16164
rect 23431 16133 23443 16136
rect 23385 16127 23443 16133
rect 23842 16124 23848 16136
rect 23900 16164 23906 16176
rect 24394 16164 24400 16176
rect 23900 16136 24400 16164
rect 23900 16124 23906 16136
rect 24394 16124 24400 16136
rect 24452 16124 24458 16176
rect 25038 16124 25044 16176
rect 25096 16124 25102 16176
rect 27522 16164 27528 16176
rect 27483 16136 27528 16164
rect 27522 16124 27528 16136
rect 27580 16124 27586 16176
rect 30282 16124 30288 16176
rect 30340 16164 30346 16176
rect 31205 16167 31263 16173
rect 31205 16164 31217 16167
rect 30340 16136 31217 16164
rect 30340 16124 30346 16136
rect 31205 16133 31217 16136
rect 31251 16133 31263 16167
rect 31205 16127 31263 16133
rect 31389 16167 31447 16173
rect 31389 16133 31401 16167
rect 31435 16164 31447 16167
rect 32944 16167 33002 16173
rect 31435 16136 32628 16164
rect 31435 16133 31447 16136
rect 31389 16127 31447 16133
rect 19628 16068 20576 16096
rect 18601 16059 18659 16065
rect 20622 16056 20628 16108
rect 20680 16096 20686 16108
rect 20809 16099 20867 16105
rect 20680 16068 20725 16096
rect 20680 16056 20686 16068
rect 20809 16065 20821 16099
rect 20855 16065 20867 16099
rect 20809 16059 20867 16065
rect 20824 16028 20852 16059
rect 22462 16056 22468 16108
rect 22520 16096 22526 16108
rect 22557 16099 22615 16105
rect 22557 16096 22569 16099
rect 22520 16068 22569 16096
rect 22520 16056 22526 16068
rect 22557 16065 22569 16068
rect 22603 16065 22615 16099
rect 22557 16059 22615 16065
rect 22741 16099 22799 16105
rect 22741 16065 22753 16099
rect 22787 16065 22799 16099
rect 22741 16059 22799 16065
rect 24121 16099 24179 16105
rect 24121 16065 24133 16099
rect 24167 16096 24179 16099
rect 25056 16096 25084 16124
rect 24167 16068 25084 16096
rect 25308 16099 25366 16105
rect 24167 16065 24179 16068
rect 24121 16059 24179 16065
rect 25308 16065 25320 16099
rect 25354 16096 25366 16099
rect 26142 16096 26148 16108
rect 25354 16068 26148 16096
rect 25354 16065 25366 16068
rect 25308 16059 25366 16065
rect 21910 16028 21916 16040
rect 20824 16000 21916 16028
rect 21910 15988 21916 16000
rect 21968 16028 21974 16040
rect 22756 16028 22784 16059
rect 26142 16056 26148 16068
rect 26200 16056 26206 16108
rect 27062 16056 27068 16108
rect 27120 16096 27126 16108
rect 27157 16099 27215 16105
rect 27157 16096 27169 16099
rect 27120 16068 27169 16096
rect 27120 16056 27126 16068
rect 27157 16065 27169 16068
rect 27203 16065 27215 16099
rect 27157 16059 27215 16065
rect 27985 16099 28043 16105
rect 27985 16065 27997 16099
rect 28031 16096 28043 16099
rect 28350 16096 28356 16108
rect 28031 16068 28356 16096
rect 28031 16065 28043 16068
rect 27985 16059 28043 16065
rect 21968 16000 22784 16028
rect 21968 15988 21974 16000
rect 24854 15988 24860 16040
rect 24912 16028 24918 16040
rect 25041 16031 25099 16037
rect 25041 16028 25053 16031
rect 24912 16000 25053 16028
rect 24912 15988 24918 16000
rect 25041 15997 25053 16000
rect 25087 15997 25099 16031
rect 26973 16031 27031 16037
rect 26973 16028 26985 16031
rect 25041 15991 25099 15997
rect 26436 16000 26985 16028
rect 18141 15963 18199 15969
rect 18141 15929 18153 15963
rect 18187 15929 18199 15963
rect 18141 15923 18199 15929
rect 20070 15920 20076 15972
rect 20128 15960 20134 15972
rect 20898 15960 20904 15972
rect 20128 15932 20904 15960
rect 20128 15920 20134 15932
rect 20898 15920 20904 15932
rect 20956 15920 20962 15972
rect 22462 15920 22468 15972
rect 22520 15960 22526 15972
rect 24305 15963 24363 15969
rect 24305 15960 24317 15963
rect 22520 15932 24317 15960
rect 22520 15920 22526 15932
rect 24305 15929 24317 15932
rect 24351 15960 24363 15963
rect 24486 15960 24492 15972
rect 24351 15932 24492 15960
rect 24351 15929 24363 15932
rect 24305 15923 24363 15929
rect 24486 15920 24492 15932
rect 24544 15920 24550 15972
rect 26436 15969 26464 16000
rect 26973 15997 26985 16000
rect 27019 15997 27031 16031
rect 27172 16028 27200 16059
rect 28350 16056 28356 16068
rect 28408 16056 28414 16108
rect 28442 16056 28448 16108
rect 28500 16096 28506 16108
rect 28721 16099 28779 16105
rect 28721 16096 28733 16099
rect 28500 16068 28733 16096
rect 28500 16056 28506 16068
rect 28721 16065 28733 16068
rect 28767 16065 28779 16099
rect 28902 16096 28908 16108
rect 28863 16068 28908 16096
rect 28721 16059 28779 16065
rect 28902 16056 28908 16068
rect 28960 16056 28966 16108
rect 30377 16099 30435 16105
rect 30377 16065 30389 16099
rect 30423 16065 30435 16099
rect 30377 16059 30435 16065
rect 30561 16099 30619 16105
rect 30561 16065 30573 16099
rect 30607 16096 30619 16099
rect 31220 16096 31248 16127
rect 32398 16096 32404 16108
rect 30607 16068 31156 16096
rect 31220 16068 32404 16096
rect 30607 16065 30619 16068
rect 30561 16059 30619 16065
rect 28077 16031 28135 16037
rect 28077 16028 28089 16031
rect 27172 16000 28089 16028
rect 26973 15991 27031 15997
rect 27908 15972 27936 16000
rect 28077 15997 28089 16000
rect 28123 16028 28135 16031
rect 28166 16028 28172 16040
rect 28123 16000 28172 16028
rect 28123 15997 28135 16000
rect 28077 15991 28135 15997
rect 28166 15988 28172 16000
rect 28224 15988 28230 16040
rect 28261 16031 28319 16037
rect 28261 15997 28273 16031
rect 28307 16028 28319 16031
rect 28534 16028 28540 16040
rect 28307 16000 28540 16028
rect 28307 15997 28319 16000
rect 28261 15991 28319 15997
rect 28534 15988 28540 16000
rect 28592 15988 28598 16040
rect 30392 16028 30420 16059
rect 30926 16028 30932 16040
rect 30392 16000 30932 16028
rect 30926 15988 30932 16000
rect 30984 15988 30990 16040
rect 26421 15963 26479 15969
rect 26421 15929 26433 15963
rect 26467 15929 26479 15963
rect 26421 15923 26479 15929
rect 27890 15920 27896 15972
rect 27948 15920 27954 15972
rect 31128 15960 31156 16068
rect 32398 16056 32404 16068
rect 32456 16056 32462 16108
rect 32306 15960 32312 15972
rect 31128 15932 32312 15960
rect 32306 15920 32312 15932
rect 32364 15920 32370 15972
rect 15286 15892 15292 15904
rect 14292 15864 15292 15892
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 20717 15895 20775 15901
rect 20717 15861 20729 15895
rect 20763 15892 20775 15895
rect 21082 15892 21088 15904
rect 20763 15864 21088 15892
rect 20763 15861 20775 15864
rect 20717 15855 20775 15861
rect 21082 15852 21088 15864
rect 21140 15852 21146 15904
rect 22554 15892 22560 15904
rect 22515 15864 22560 15892
rect 22554 15852 22560 15864
rect 22612 15852 22618 15904
rect 23474 15852 23480 15904
rect 23532 15892 23538 15904
rect 23569 15895 23627 15901
rect 23569 15892 23581 15895
rect 23532 15864 23581 15892
rect 23532 15852 23538 15864
rect 23569 15861 23581 15864
rect 23615 15861 23627 15895
rect 23569 15855 23627 15861
rect 27433 15895 27491 15901
rect 27433 15861 27445 15895
rect 27479 15892 27491 15895
rect 27706 15892 27712 15904
rect 27479 15864 27712 15892
rect 27479 15861 27491 15864
rect 27433 15855 27491 15861
rect 27706 15852 27712 15864
rect 27764 15852 27770 15904
rect 28166 15852 28172 15904
rect 28224 15892 28230 15904
rect 30742 15892 30748 15904
rect 28224 15864 28269 15892
rect 30703 15864 30748 15892
rect 28224 15852 28230 15864
rect 30742 15852 30748 15864
rect 30800 15852 30806 15904
rect 31573 15895 31631 15901
rect 31573 15861 31585 15895
rect 31619 15892 31631 15895
rect 32490 15892 32496 15904
rect 31619 15864 32496 15892
rect 31619 15861 31631 15864
rect 31573 15855 31631 15861
rect 32490 15852 32496 15864
rect 32548 15852 32554 15904
rect 32600 15892 32628 16136
rect 32944 16133 32956 16167
rect 32990 16164 33002 16167
rect 34532 16164 34560 16204
rect 36357 16201 36369 16204
rect 36403 16201 36415 16235
rect 36357 16195 36415 16201
rect 32990 16136 34560 16164
rect 32990 16133 33002 16136
rect 32944 16127 33002 16133
rect 34422 16096 34428 16108
rect 32692 16068 34428 16096
rect 32692 16040 32720 16068
rect 34422 16056 34428 16068
rect 34480 16096 34486 16108
rect 34517 16099 34575 16105
rect 34517 16096 34529 16099
rect 34480 16068 34529 16096
rect 34480 16056 34486 16068
rect 34517 16065 34529 16068
rect 34563 16065 34575 16099
rect 34517 16059 34575 16065
rect 34606 16056 34612 16108
rect 34664 16096 34670 16108
rect 34773 16099 34831 16105
rect 34773 16096 34785 16099
rect 34664 16068 34785 16096
rect 34664 16056 34670 16068
rect 34773 16065 34785 16068
rect 34819 16065 34831 16099
rect 34773 16059 34831 16065
rect 36446 16056 36452 16108
rect 36504 16096 36510 16108
rect 36541 16099 36599 16105
rect 36541 16096 36553 16099
rect 36504 16068 36553 16096
rect 36504 16056 36510 16068
rect 36541 16065 36553 16068
rect 36587 16065 36599 16099
rect 36541 16059 36599 16065
rect 32674 15988 32680 16040
rect 32732 16028 32738 16040
rect 32732 16000 32777 16028
rect 32732 15988 32738 16000
rect 33686 15920 33692 15972
rect 33744 15960 33750 15972
rect 33744 15932 34560 15960
rect 33744 15920 33750 15932
rect 34238 15892 34244 15904
rect 32600 15864 34244 15892
rect 34238 15852 34244 15864
rect 34296 15852 34302 15904
rect 34532 15892 34560 15932
rect 35710 15892 35716 15904
rect 34532 15864 35716 15892
rect 35710 15852 35716 15864
rect 35768 15852 35774 15904
rect 35894 15892 35900 15904
rect 35855 15864 35900 15892
rect 35894 15852 35900 15864
rect 35952 15852 35958 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 3237 15691 3295 15697
rect 3237 15657 3249 15691
rect 3283 15688 3295 15691
rect 3283 15660 7696 15688
rect 3283 15657 3295 15660
rect 3237 15651 3295 15657
rect 1854 15552 1860 15564
rect 1815 15524 1860 15552
rect 1854 15512 1860 15524
rect 1912 15512 1918 15564
rect 6730 15512 6736 15564
rect 6788 15552 6794 15564
rect 6788 15524 7512 15552
rect 6788 15512 6794 15524
rect 3786 15484 3792 15496
rect 3699 15456 3792 15484
rect 3786 15444 3792 15456
rect 3844 15484 3850 15496
rect 5629 15487 5687 15493
rect 5629 15484 5641 15487
rect 3844 15456 5641 15484
rect 3844 15444 3850 15456
rect 5629 15453 5641 15456
rect 5675 15484 5687 15487
rect 6822 15484 6828 15496
rect 5675 15456 6828 15484
rect 5675 15453 5687 15456
rect 5629 15447 5687 15453
rect 6822 15444 6828 15456
rect 6880 15444 6886 15496
rect 2124 15419 2182 15425
rect 2124 15385 2136 15419
rect 2170 15416 2182 15419
rect 3878 15416 3884 15428
rect 2170 15388 3884 15416
rect 2170 15385 2182 15388
rect 2124 15379 2182 15385
rect 3878 15376 3884 15388
rect 3936 15376 3942 15428
rect 4056 15419 4114 15425
rect 4056 15385 4068 15419
rect 4102 15416 4114 15419
rect 4798 15416 4804 15428
rect 4102 15388 4804 15416
rect 4102 15385 4114 15388
rect 4056 15379 4114 15385
rect 4798 15376 4804 15388
rect 4856 15376 4862 15428
rect 5902 15425 5908 15428
rect 5896 15416 5908 15425
rect 5863 15388 5908 15416
rect 5896 15379 5908 15388
rect 5902 15376 5908 15379
rect 5960 15376 5966 15428
rect 5994 15376 6000 15428
rect 6052 15416 6058 15428
rect 7484 15425 7512 15524
rect 7668 15493 7696 15660
rect 9766 15648 9772 15700
rect 9824 15688 9830 15700
rect 10870 15688 10876 15700
rect 9824 15660 10876 15688
rect 9824 15648 9830 15660
rect 10870 15648 10876 15660
rect 10928 15688 10934 15700
rect 11146 15688 11152 15700
rect 10928 15660 11152 15688
rect 10928 15648 10934 15660
rect 11146 15648 11152 15660
rect 11204 15648 11210 15700
rect 12710 15688 12716 15700
rect 12671 15660 12716 15688
rect 12710 15648 12716 15660
rect 12768 15648 12774 15700
rect 14921 15691 14979 15697
rect 14921 15657 14933 15691
rect 14967 15688 14979 15691
rect 15102 15688 15108 15700
rect 14967 15660 15108 15688
rect 14967 15657 14979 15660
rect 14921 15651 14979 15657
rect 15102 15648 15108 15660
rect 15160 15648 15166 15700
rect 15378 15648 15384 15700
rect 15436 15688 15442 15700
rect 15473 15691 15531 15697
rect 15473 15688 15485 15691
rect 15436 15660 15485 15688
rect 15436 15648 15442 15660
rect 15473 15657 15485 15660
rect 15519 15657 15531 15691
rect 15473 15651 15531 15657
rect 17681 15691 17739 15697
rect 17681 15657 17693 15691
rect 17727 15688 17739 15691
rect 18138 15688 18144 15700
rect 17727 15660 18144 15688
rect 17727 15657 17739 15660
rect 17681 15651 17739 15657
rect 18138 15648 18144 15660
rect 18196 15648 18202 15700
rect 18598 15648 18604 15700
rect 18656 15688 18662 15700
rect 19797 15691 19855 15697
rect 19797 15688 19809 15691
rect 18656 15660 19809 15688
rect 18656 15648 18662 15660
rect 19797 15657 19809 15660
rect 19843 15688 19855 15691
rect 20622 15688 20628 15700
rect 19843 15660 20628 15688
rect 19843 15657 19855 15660
rect 19797 15651 19855 15657
rect 20622 15648 20628 15660
rect 20680 15648 20686 15700
rect 23290 15688 23296 15700
rect 23251 15660 23296 15688
rect 23290 15648 23296 15660
rect 23348 15648 23354 15700
rect 26142 15688 26148 15700
rect 26103 15660 26148 15688
rect 26142 15648 26148 15660
rect 26200 15648 26206 15700
rect 27614 15688 27620 15700
rect 27575 15660 27620 15688
rect 27614 15648 27620 15660
rect 27672 15648 27678 15700
rect 36081 15691 36139 15697
rect 36081 15688 36093 15691
rect 32140 15660 36093 15688
rect 10778 15580 10784 15632
rect 10836 15620 10842 15632
rect 11238 15620 11244 15632
rect 10836 15592 11244 15620
rect 10836 15580 10842 15592
rect 11238 15580 11244 15592
rect 11296 15620 11302 15632
rect 11977 15623 12035 15629
rect 11977 15620 11989 15623
rect 11296 15592 11989 15620
rect 11296 15580 11302 15592
rect 11977 15589 11989 15592
rect 12023 15589 12035 15623
rect 22462 15620 22468 15632
rect 11977 15583 12035 15589
rect 17696 15592 22468 15620
rect 13262 15552 13268 15564
rect 13096 15524 13268 15552
rect 7653 15487 7711 15493
rect 7653 15453 7665 15487
rect 7699 15453 7711 15487
rect 7653 15447 7711 15453
rect 8938 15444 8944 15496
rect 8996 15484 9002 15496
rect 9125 15487 9183 15493
rect 9125 15484 9137 15487
rect 8996 15456 9137 15484
rect 8996 15444 9002 15456
rect 9125 15453 9137 15456
rect 9171 15453 9183 15487
rect 9766 15484 9772 15496
rect 9727 15456 9772 15484
rect 9125 15447 9183 15453
rect 9766 15444 9772 15456
rect 9824 15444 9830 15496
rect 10036 15487 10094 15493
rect 10036 15453 10048 15487
rect 10082 15484 10094 15487
rect 10318 15484 10324 15496
rect 10082 15456 10324 15484
rect 10082 15453 10094 15456
rect 10036 15447 10094 15453
rect 10318 15444 10324 15456
rect 10376 15444 10382 15496
rect 10502 15444 10508 15496
rect 10560 15484 10566 15496
rect 12066 15484 12072 15496
rect 10560 15456 12072 15484
rect 10560 15444 10566 15456
rect 12066 15444 12072 15456
rect 12124 15484 12130 15496
rect 12894 15484 12900 15496
rect 12124 15456 12900 15484
rect 12124 15444 12130 15456
rect 12894 15444 12900 15456
rect 12952 15484 12958 15496
rect 13096 15493 13124 15524
rect 13262 15512 13268 15524
rect 13320 15552 13326 15564
rect 14090 15552 14096 15564
rect 13320 15524 14096 15552
rect 13320 15512 13326 15524
rect 14090 15512 14096 15524
rect 14148 15512 14154 15564
rect 15028 15524 15700 15552
rect 12989 15487 13047 15493
rect 12989 15484 13001 15487
rect 12952 15456 13001 15484
rect 12952 15444 12958 15456
rect 12989 15453 13001 15456
rect 13035 15453 13047 15487
rect 12989 15447 13047 15453
rect 13081 15487 13139 15493
rect 13081 15453 13093 15487
rect 13127 15453 13139 15487
rect 13081 15447 13139 15453
rect 13170 15444 13176 15496
rect 13228 15484 13234 15496
rect 13357 15487 13415 15493
rect 13228 15456 13273 15484
rect 13228 15444 13234 15456
rect 13357 15453 13369 15487
rect 13403 15453 13415 15487
rect 13357 15447 13415 15453
rect 14829 15487 14887 15493
rect 14829 15453 14841 15487
rect 14875 15484 14887 15487
rect 14918 15484 14924 15496
rect 14875 15456 14924 15484
rect 14875 15453 14887 15456
rect 14829 15447 14887 15453
rect 7469 15419 7527 15425
rect 6052 15388 7144 15416
rect 6052 15376 6058 15388
rect 5169 15351 5227 15357
rect 5169 15317 5181 15351
rect 5215 15348 5227 15351
rect 6546 15348 6552 15360
rect 5215 15320 6552 15348
rect 5215 15317 5227 15320
rect 5169 15311 5227 15317
rect 6546 15308 6552 15320
rect 6604 15308 6610 15360
rect 7006 15348 7012 15360
rect 6967 15320 7012 15348
rect 7006 15308 7012 15320
rect 7064 15308 7070 15360
rect 7116 15348 7144 15388
rect 7469 15385 7481 15419
rect 7515 15416 7527 15419
rect 11606 15416 11612 15428
rect 7515 15388 8892 15416
rect 11567 15388 11612 15416
rect 7515 15385 7527 15388
rect 7469 15379 7527 15385
rect 8864 15360 8892 15388
rect 11606 15376 11612 15388
rect 11664 15376 11670 15428
rect 11793 15419 11851 15425
rect 11793 15385 11805 15419
rect 11839 15385 11851 15419
rect 11793 15379 11851 15385
rect 7837 15351 7895 15357
rect 7837 15348 7849 15351
rect 7116 15320 7849 15348
rect 7837 15317 7849 15320
rect 7883 15317 7895 15351
rect 7837 15311 7895 15317
rect 8846 15308 8852 15360
rect 8904 15348 8910 15360
rect 8941 15351 8999 15357
rect 8941 15348 8953 15351
rect 8904 15320 8953 15348
rect 8904 15308 8910 15320
rect 8941 15317 8953 15320
rect 8987 15317 8999 15351
rect 8941 15311 8999 15317
rect 11149 15351 11207 15357
rect 11149 15317 11161 15351
rect 11195 15348 11207 15351
rect 11808 15348 11836 15379
rect 12710 15376 12716 15428
rect 12768 15416 12774 15428
rect 13372 15416 13400 15447
rect 14918 15444 14924 15456
rect 14976 15444 14982 15496
rect 15028 15493 15056 15524
rect 15672 15493 15700 15524
rect 15013 15487 15071 15493
rect 15013 15453 15025 15487
rect 15059 15453 15071 15487
rect 15013 15447 15071 15453
rect 15473 15487 15531 15493
rect 15473 15453 15485 15487
rect 15519 15453 15531 15487
rect 15473 15447 15531 15453
rect 15657 15487 15715 15493
rect 15657 15453 15669 15487
rect 15703 15484 15715 15487
rect 16022 15484 16028 15496
rect 15703 15456 16028 15484
rect 15703 15453 15715 15456
rect 15657 15447 15715 15453
rect 12768 15388 13400 15416
rect 15488 15416 15516 15447
rect 16022 15444 16028 15456
rect 16080 15444 16086 15496
rect 17696 15493 17724 15592
rect 22462 15580 22468 15592
rect 22520 15580 22526 15632
rect 31481 15623 31539 15629
rect 31481 15589 31493 15623
rect 31527 15620 31539 15623
rect 31938 15620 31944 15632
rect 31527 15592 31944 15620
rect 31527 15589 31539 15592
rect 31481 15583 31539 15589
rect 31938 15580 31944 15592
rect 31996 15580 32002 15632
rect 20438 15512 20444 15564
rect 20496 15552 20502 15564
rect 22554 15552 22560 15564
rect 20496 15524 21956 15552
rect 20496 15512 20502 15524
rect 17681 15487 17739 15493
rect 17681 15453 17693 15487
rect 17727 15453 17739 15487
rect 17862 15484 17868 15496
rect 17823 15456 17868 15484
rect 17681 15447 17739 15453
rect 17862 15444 17868 15456
rect 17920 15444 17926 15496
rect 21008 15493 21036 15524
rect 20901 15487 20959 15493
rect 20901 15484 20913 15487
rect 19306 15456 20913 15484
rect 17954 15416 17960 15428
rect 15488 15388 17960 15416
rect 12768 15376 12774 15388
rect 17954 15376 17960 15388
rect 18012 15376 18018 15428
rect 11195 15320 11836 15348
rect 11195 15317 11207 15320
rect 11149 15311 11207 15317
rect 12894 15308 12900 15360
rect 12952 15348 12958 15360
rect 16758 15348 16764 15360
rect 12952 15320 16764 15348
rect 12952 15308 12958 15320
rect 16758 15308 16764 15320
rect 16816 15348 16822 15360
rect 19306 15348 19334 15456
rect 20901 15453 20913 15456
rect 20947 15453 20959 15487
rect 20901 15447 20959 15453
rect 20993 15487 21051 15493
rect 20993 15453 21005 15487
rect 21039 15453 21051 15487
rect 20993 15447 21051 15453
rect 21082 15444 21088 15496
rect 21140 15484 21146 15496
rect 21140 15456 21185 15484
rect 21140 15444 21146 15456
rect 21266 15444 21272 15496
rect 21324 15484 21330 15496
rect 21928 15493 21956 15524
rect 22204 15524 22560 15552
rect 21913 15487 21971 15493
rect 21324 15456 21369 15484
rect 21324 15444 21330 15456
rect 21913 15453 21925 15487
rect 21959 15453 21971 15487
rect 21913 15447 21971 15453
rect 22002 15444 22008 15496
rect 22060 15484 22066 15496
rect 22204 15493 22232 15524
rect 22554 15512 22560 15524
rect 22612 15512 22618 15564
rect 30834 15552 30840 15564
rect 30484 15524 30840 15552
rect 22189 15487 22247 15493
rect 22060 15456 22105 15484
rect 22060 15444 22066 15456
rect 22189 15453 22201 15487
rect 22235 15453 22247 15487
rect 22189 15447 22247 15453
rect 22281 15487 22339 15493
rect 22281 15453 22293 15487
rect 22327 15453 22339 15487
rect 23474 15484 23480 15496
rect 23435 15456 23480 15484
rect 22281 15447 22339 15453
rect 19702 15416 19708 15428
rect 19663 15388 19708 15416
rect 19702 15376 19708 15388
rect 19760 15376 19766 15428
rect 22296 15416 22324 15447
rect 23474 15444 23480 15456
rect 23532 15444 23538 15496
rect 24670 15444 24676 15496
rect 24728 15484 24734 15496
rect 24857 15487 24915 15493
rect 24857 15484 24869 15487
rect 24728 15456 24869 15484
rect 24728 15444 24734 15456
rect 24857 15453 24869 15456
rect 24903 15453 24915 15487
rect 26142 15484 26148 15496
rect 26103 15456 26148 15484
rect 24857 15447 24915 15453
rect 26142 15444 26148 15456
rect 26200 15444 26206 15496
rect 26329 15487 26387 15493
rect 26329 15453 26341 15487
rect 26375 15484 26387 15487
rect 27522 15484 27528 15496
rect 26375 15456 27528 15484
rect 26375 15453 26387 15456
rect 26329 15447 26387 15453
rect 27522 15444 27528 15456
rect 27580 15444 27586 15496
rect 27617 15487 27675 15493
rect 27617 15453 27629 15487
rect 27663 15453 27675 15487
rect 27617 15447 27675 15453
rect 27801 15487 27859 15493
rect 27801 15453 27813 15487
rect 27847 15484 27859 15487
rect 28166 15484 28172 15496
rect 27847 15456 28172 15484
rect 27847 15453 27859 15456
rect 27801 15447 27859 15453
rect 24688 15416 24716 15444
rect 27632 15416 27660 15447
rect 28166 15444 28172 15456
rect 28224 15484 28230 15496
rect 28810 15484 28816 15496
rect 28224 15456 28816 15484
rect 28224 15444 28230 15456
rect 28810 15444 28816 15456
rect 28868 15444 28874 15496
rect 29825 15487 29883 15493
rect 29825 15453 29837 15487
rect 29871 15453 29883 15487
rect 30282 15484 30288 15496
rect 30243 15456 30288 15484
rect 29825 15447 29883 15453
rect 22296 15388 24716 15416
rect 26988 15388 27660 15416
rect 29840 15416 29868 15447
rect 30282 15444 30288 15456
rect 30340 15444 30346 15496
rect 30484 15493 30512 15524
rect 30834 15512 30840 15524
rect 30892 15512 30898 15564
rect 31846 15552 31852 15564
rect 31036 15524 31852 15552
rect 30469 15487 30527 15493
rect 30469 15453 30481 15487
rect 30515 15453 30527 15487
rect 30469 15447 30527 15453
rect 30653 15487 30711 15493
rect 30653 15453 30665 15487
rect 30699 15484 30711 15487
rect 31036 15484 31064 15524
rect 31846 15512 31852 15524
rect 31904 15512 31910 15564
rect 31588 15484 31754 15494
rect 32140 15493 32168 15660
rect 36081 15657 36093 15660
rect 36127 15657 36139 15691
rect 36081 15651 36139 15657
rect 33870 15580 33876 15632
rect 33928 15620 33934 15632
rect 34149 15623 34207 15629
rect 34149 15620 34161 15623
rect 33928 15592 34161 15620
rect 33928 15580 33934 15592
rect 34149 15589 34161 15592
rect 34195 15589 34207 15623
rect 34149 15583 34207 15589
rect 36538 15552 36544 15564
rect 36499 15524 36544 15552
rect 36538 15512 36544 15524
rect 36596 15512 36602 15564
rect 32125 15487 32183 15493
rect 30699 15456 31064 15484
rect 31128 15466 31984 15484
rect 31128 15456 31616 15466
rect 31726 15456 31984 15466
rect 30699 15453 30711 15456
rect 30653 15447 30711 15453
rect 30834 15416 30840 15428
rect 29840 15388 30840 15416
rect 26988 15360 27016 15388
rect 30834 15376 30840 15388
rect 30892 15376 30898 15428
rect 31128 15425 31156 15456
rect 31113 15419 31171 15425
rect 31113 15385 31125 15419
rect 31159 15385 31171 15419
rect 31113 15379 31171 15385
rect 31297 15419 31355 15425
rect 31297 15385 31309 15419
rect 31343 15416 31355 15419
rect 31846 15416 31852 15428
rect 31343 15388 31852 15416
rect 31343 15385 31355 15388
rect 31297 15379 31355 15385
rect 31846 15376 31852 15388
rect 31904 15376 31910 15428
rect 31956 15425 31984 15456
rect 32125 15453 32137 15487
rect 32171 15453 32183 15487
rect 32125 15447 32183 15453
rect 32674 15444 32680 15496
rect 32732 15484 32738 15496
rect 32769 15487 32827 15493
rect 32769 15484 32781 15487
rect 32732 15456 32781 15484
rect 32732 15444 32738 15456
rect 32769 15453 32781 15456
rect 32815 15453 32827 15487
rect 32769 15447 32827 15453
rect 33036 15487 33094 15493
rect 33036 15453 33048 15487
rect 33082 15484 33094 15487
rect 33082 15456 33180 15484
rect 33082 15453 33094 15456
rect 33036 15447 33094 15453
rect 31941 15419 31999 15425
rect 31941 15385 31953 15419
rect 31987 15385 31999 15419
rect 31941 15379 31999 15385
rect 16816 15320 19334 15348
rect 20625 15351 20683 15357
rect 16816 15308 16822 15320
rect 20625 15317 20637 15351
rect 20671 15348 20683 15351
rect 20714 15348 20720 15360
rect 20671 15320 20720 15348
rect 20671 15317 20683 15320
rect 20625 15311 20683 15317
rect 20714 15308 20720 15320
rect 20772 15308 20778 15360
rect 21729 15351 21787 15357
rect 21729 15317 21741 15351
rect 21775 15348 21787 15351
rect 22094 15348 22100 15360
rect 21775 15320 22100 15348
rect 21775 15317 21787 15320
rect 21729 15311 21787 15317
rect 22094 15308 22100 15320
rect 22152 15308 22158 15360
rect 24949 15351 25007 15357
rect 24949 15317 24961 15351
rect 24995 15348 25007 15351
rect 25038 15348 25044 15360
rect 24995 15320 25044 15348
rect 24995 15317 25007 15320
rect 24949 15311 25007 15317
rect 25038 15308 25044 15320
rect 25096 15348 25102 15360
rect 26970 15348 26976 15360
rect 25096 15320 26976 15348
rect 25096 15308 25102 15320
rect 26970 15308 26976 15320
rect 27028 15308 27034 15360
rect 29641 15351 29699 15357
rect 29641 15317 29653 15351
rect 29687 15348 29699 15351
rect 31754 15348 31760 15360
rect 29687 15320 31760 15348
rect 29687 15317 29699 15320
rect 29641 15311 29699 15317
rect 31754 15308 31760 15320
rect 31812 15308 31818 15360
rect 31956 15348 31984 15379
rect 32122 15348 32128 15360
rect 31956 15320 32128 15348
rect 32122 15308 32128 15320
rect 32180 15308 32186 15360
rect 32309 15351 32367 15357
rect 32309 15317 32321 15351
rect 32355 15348 32367 15351
rect 32858 15348 32864 15360
rect 32355 15320 32864 15348
rect 32355 15317 32367 15320
rect 32309 15311 32367 15317
rect 32858 15308 32864 15320
rect 32916 15308 32922 15360
rect 33152 15348 33180 15456
rect 34422 15444 34428 15496
rect 34480 15484 34486 15496
rect 34701 15487 34759 15493
rect 34701 15484 34713 15487
rect 34480 15456 34713 15484
rect 34480 15444 34486 15456
rect 34701 15453 34713 15456
rect 34747 15453 34759 15487
rect 34701 15447 34759 15453
rect 34238 15376 34244 15428
rect 34296 15416 34302 15428
rect 34946 15419 35004 15425
rect 34946 15416 34958 15419
rect 34296 15388 34958 15416
rect 34296 15376 34302 15388
rect 34946 15385 34958 15388
rect 34992 15385 35004 15419
rect 34946 15379 35004 15385
rect 35986 15376 35992 15428
rect 36044 15416 36050 15428
rect 36786 15419 36844 15425
rect 36786 15416 36798 15419
rect 36044 15388 36798 15416
rect 36044 15376 36050 15388
rect 36786 15385 36798 15388
rect 36832 15385 36844 15419
rect 36786 15379 36844 15385
rect 33778 15348 33784 15360
rect 33152 15320 33784 15348
rect 33778 15308 33784 15320
rect 33836 15308 33842 15360
rect 34514 15308 34520 15360
rect 34572 15348 34578 15360
rect 37921 15351 37979 15357
rect 37921 15348 37933 15351
rect 34572 15320 37933 15348
rect 34572 15308 34578 15320
rect 37921 15317 37933 15320
rect 37967 15317 37979 15351
rect 37921 15311 37979 15317
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 3878 15104 3884 15156
rect 3936 15144 3942 15156
rect 4801 15147 4859 15153
rect 4801 15144 4813 15147
rect 3936 15116 4813 15144
rect 3936 15104 3942 15116
rect 4801 15113 4813 15116
rect 4847 15113 4859 15147
rect 6733 15147 6791 15153
rect 4801 15107 4859 15113
rect 4908 15116 6132 15144
rect 2952 15079 3010 15085
rect 2952 15045 2964 15079
rect 2998 15076 3010 15079
rect 4908 15076 4936 15116
rect 5994 15076 6000 15088
rect 2998 15048 4936 15076
rect 5000 15048 6000 15076
rect 2998 15045 3010 15048
rect 2952 15039 3010 15045
rect 2682 15008 2688 15020
rect 2643 14980 2688 15008
rect 2682 14968 2688 14980
rect 2740 14968 2746 15020
rect 5000 15017 5028 15048
rect 5994 15036 6000 15048
rect 6052 15036 6058 15088
rect 6104 15076 6132 15116
rect 6733 15113 6745 15147
rect 6779 15144 6791 15147
rect 7374 15144 7380 15156
rect 6779 15116 7380 15144
rect 6779 15113 6791 15116
rect 6733 15107 6791 15113
rect 7374 15104 7380 15116
rect 7432 15104 7438 15156
rect 8018 15144 8024 15156
rect 7979 15116 8024 15144
rect 8018 15104 8024 15116
rect 8076 15104 8082 15156
rect 8202 15104 8208 15156
rect 8260 15104 8266 15156
rect 13262 15104 13268 15156
rect 13320 15144 13326 15156
rect 13357 15147 13415 15153
rect 13357 15144 13369 15147
rect 13320 15116 13369 15144
rect 13320 15104 13326 15116
rect 13357 15113 13369 15116
rect 13403 15113 13415 15147
rect 17589 15147 17647 15153
rect 17589 15144 17601 15147
rect 13357 15107 13415 15113
rect 15120 15116 17601 15144
rect 6914 15076 6920 15088
rect 6104 15048 6920 15076
rect 6914 15036 6920 15048
rect 6972 15036 6978 15088
rect 7193 15079 7251 15085
rect 7193 15045 7205 15079
rect 7239 15076 7251 15079
rect 8220 15076 8248 15104
rect 7239 15048 8248 15076
rect 8956 15048 10180 15076
rect 7239 15045 7251 15048
rect 7193 15039 7251 15045
rect 8956 15020 8984 15048
rect 4985 15011 5043 15017
rect 4985 14977 4997 15011
rect 5031 14977 5043 15011
rect 4985 14971 5043 14977
rect 5350 14968 5356 15020
rect 5408 15008 5414 15020
rect 5445 15011 5503 15017
rect 5445 15008 5457 15011
rect 5408 14980 5457 15008
rect 5408 14968 5414 14980
rect 5445 14977 5457 14980
rect 5491 14977 5503 15011
rect 5445 14971 5503 14977
rect 5534 14968 5540 15020
rect 5592 15008 5598 15020
rect 5629 15011 5687 15017
rect 5629 15008 5641 15011
rect 5592 14980 5641 15008
rect 5592 14968 5598 14980
rect 5629 14977 5641 14980
rect 5675 14977 5687 15011
rect 6362 15008 6368 15020
rect 6323 14980 6368 15008
rect 5629 14971 5687 14977
rect 6362 14968 6368 14980
rect 6420 14968 6426 15020
rect 6549 15011 6607 15017
rect 6549 14977 6561 15011
rect 6595 14977 6607 15011
rect 6549 14971 6607 14977
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 14977 7435 15011
rect 7377 14971 7435 14977
rect 6564 14940 6592 14971
rect 4080 14912 6592 14940
rect 4080 14881 4108 14912
rect 6638 14900 6644 14952
rect 6696 14940 6702 14952
rect 7392 14940 7420 14971
rect 7834 14968 7840 15020
rect 7892 15008 7898 15020
rect 8205 15011 8263 15017
rect 8205 15008 8217 15011
rect 7892 14980 8217 15008
rect 7892 14968 7898 14980
rect 8205 14977 8217 14980
rect 8251 14977 8263 15011
rect 8205 14971 8263 14977
rect 8849 15011 8907 15017
rect 8849 14977 8861 15011
rect 8895 15008 8907 15011
rect 8938 15008 8944 15020
rect 8895 14980 8944 15008
rect 8895 14977 8907 14980
rect 8849 14971 8907 14977
rect 8938 14968 8944 14980
rect 8996 14968 9002 15020
rect 9030 14968 9036 15020
rect 9088 15008 9094 15020
rect 10152 15017 10180 15048
rect 11606 15036 11612 15088
rect 11664 15076 11670 15088
rect 12989 15079 13047 15085
rect 12989 15076 13001 15079
rect 11664 15048 13001 15076
rect 11664 15036 11670 15048
rect 12989 15045 13001 15048
rect 13035 15045 13047 15079
rect 12989 15039 13047 15045
rect 13173 15079 13231 15085
rect 13173 15045 13185 15079
rect 13219 15076 13231 15079
rect 13538 15076 13544 15088
rect 13219 15048 13544 15076
rect 13219 15045 13231 15048
rect 13173 15039 13231 15045
rect 13538 15036 13544 15048
rect 13596 15036 13602 15088
rect 9493 15011 9551 15017
rect 9493 15008 9505 15011
rect 9088 14980 9505 15008
rect 9088 14968 9094 14980
rect 9493 14977 9505 14980
rect 9539 14977 9551 15011
rect 9493 14971 9551 14977
rect 10137 15011 10195 15017
rect 10137 14977 10149 15011
rect 10183 14977 10195 15011
rect 10137 14971 10195 14977
rect 11790 14968 11796 15020
rect 11848 15008 11854 15020
rect 15120 15008 15148 15116
rect 17589 15113 17601 15116
rect 17635 15144 17647 15147
rect 20990 15144 20996 15156
rect 17635 15116 20996 15144
rect 17635 15113 17647 15116
rect 17589 15107 17647 15113
rect 20990 15104 20996 15116
rect 21048 15104 21054 15156
rect 21266 15104 21272 15156
rect 21324 15144 21330 15156
rect 21324 15116 23612 15144
rect 21324 15104 21330 15116
rect 15197 15079 15255 15085
rect 15197 15045 15209 15079
rect 15243 15076 15255 15079
rect 16666 15076 16672 15088
rect 15243 15048 16672 15076
rect 15243 15045 15255 15048
rect 15197 15039 15255 15045
rect 16666 15036 16672 15048
rect 16724 15076 16730 15088
rect 16945 15079 17003 15085
rect 16945 15076 16957 15079
rect 16724 15048 16957 15076
rect 16724 15036 16730 15048
rect 16945 15045 16957 15048
rect 16991 15076 17003 15079
rect 18509 15079 18567 15085
rect 18509 15076 18521 15079
rect 16991 15048 18521 15076
rect 16991 15045 17003 15048
rect 16945 15039 17003 15045
rect 18509 15045 18521 15048
rect 18555 15045 18567 15079
rect 20162 15076 20168 15088
rect 18509 15039 18567 15045
rect 19260 15048 20168 15076
rect 11848 14980 15148 15008
rect 15933 15011 15991 15017
rect 11848 14968 11854 14980
rect 15933 14977 15945 15011
rect 15979 15008 15991 15011
rect 18233 15011 18291 15017
rect 15979 14980 17632 15008
rect 15979 14977 15991 14980
rect 15933 14971 15991 14977
rect 6696 14912 7420 14940
rect 6696 14900 6702 14912
rect 7926 14900 7932 14952
rect 7984 14940 7990 14952
rect 15565 14943 15623 14949
rect 7984 14912 9996 14940
rect 7984 14900 7990 14912
rect 4065 14875 4123 14881
rect 4065 14841 4077 14875
rect 4111 14841 4123 14875
rect 4065 14835 4123 14841
rect 4798 14832 4804 14884
rect 4856 14872 4862 14884
rect 9968 14881 9996 14912
rect 15565 14909 15577 14943
rect 15611 14940 15623 14943
rect 15654 14940 15660 14952
rect 15611 14912 15660 14940
rect 15611 14909 15623 14912
rect 15565 14903 15623 14909
rect 15654 14900 15660 14912
rect 15712 14900 15718 14952
rect 9309 14875 9367 14881
rect 9309 14872 9321 14875
rect 4856 14844 9321 14872
rect 4856 14832 4862 14844
rect 9309 14841 9321 14844
rect 9355 14841 9367 14875
rect 9309 14835 9367 14841
rect 9953 14875 10011 14881
rect 9953 14841 9965 14875
rect 9999 14841 10011 14875
rect 9953 14835 10011 14841
rect 10594 14832 10600 14884
rect 10652 14872 10658 14884
rect 16040 14872 16068 14980
rect 17313 14943 17371 14949
rect 17313 14909 17325 14943
rect 17359 14940 17371 14943
rect 17402 14940 17408 14952
rect 17359 14912 17408 14940
rect 17359 14909 17371 14912
rect 17313 14903 17371 14909
rect 17402 14900 17408 14912
rect 17460 14900 17466 14952
rect 17604 14940 17632 14980
rect 18233 14977 18245 15011
rect 18279 14977 18291 15011
rect 18233 14971 18291 14977
rect 17604 14912 18092 14940
rect 10652 14844 16068 14872
rect 10652 14832 10658 14844
rect 5813 14807 5871 14813
rect 5813 14773 5825 14807
rect 5859 14804 5871 14807
rect 6454 14804 6460 14816
rect 5859 14776 6460 14804
rect 5859 14773 5871 14776
rect 5813 14767 5871 14773
rect 6454 14764 6460 14776
rect 6512 14764 6518 14816
rect 6638 14764 6644 14816
rect 6696 14804 6702 14816
rect 7561 14807 7619 14813
rect 7561 14804 7573 14807
rect 6696 14776 7573 14804
rect 6696 14764 6702 14776
rect 7561 14773 7573 14776
rect 7607 14773 7619 14807
rect 7561 14767 7619 14773
rect 8202 14764 8208 14816
rect 8260 14804 8266 14816
rect 8665 14807 8723 14813
rect 8665 14804 8677 14807
rect 8260 14776 8677 14804
rect 8260 14764 8266 14776
rect 8665 14773 8677 14776
rect 8711 14773 8723 14807
rect 8665 14767 8723 14773
rect 15194 14764 15200 14816
rect 15252 14804 15258 14816
rect 15335 14807 15393 14813
rect 15335 14804 15347 14807
rect 15252 14776 15347 14804
rect 15252 14764 15258 14776
rect 15335 14773 15347 14776
rect 15381 14773 15393 14807
rect 15335 14767 15393 14773
rect 15470 14764 15476 14816
rect 15528 14804 15534 14816
rect 15528 14776 15573 14804
rect 15528 14764 15534 14776
rect 16850 14764 16856 14816
rect 16908 14804 16914 14816
rect 17083 14807 17141 14813
rect 17083 14804 17095 14807
rect 16908 14776 17095 14804
rect 16908 14764 16914 14776
rect 17083 14773 17095 14776
rect 17129 14773 17141 14807
rect 17083 14767 17141 14773
rect 17221 14807 17279 14813
rect 17221 14773 17233 14807
rect 17267 14804 17279 14807
rect 17862 14804 17868 14816
rect 17267 14776 17868 14804
rect 17267 14773 17279 14776
rect 17221 14767 17279 14773
rect 17862 14764 17868 14776
rect 17920 14764 17926 14816
rect 18064 14804 18092 14912
rect 18138 14900 18144 14952
rect 18196 14940 18202 14952
rect 18248 14940 18276 14971
rect 18322 14968 18328 15020
rect 18380 15008 18386 15020
rect 18598 15008 18604 15020
rect 18380 14980 18604 15008
rect 18380 14968 18386 14980
rect 18598 14968 18604 14980
rect 18656 14968 18662 15020
rect 19150 14940 19156 14952
rect 18196 14912 19156 14940
rect 18196 14900 18202 14912
rect 19150 14900 19156 14912
rect 19208 14900 19214 14952
rect 19260 14804 19288 15048
rect 20162 15036 20168 15048
rect 20220 15036 20226 15088
rect 22186 15076 22192 15088
rect 21836 15048 22192 15076
rect 19981 15011 20039 15017
rect 19981 14977 19993 15011
rect 20027 15008 20039 15011
rect 21266 15008 21272 15020
rect 20027 14980 21272 15008
rect 20027 14977 20039 14980
rect 19981 14971 20039 14977
rect 21266 14968 21272 14980
rect 21324 14968 21330 15020
rect 21836 15017 21864 15048
rect 22186 15036 22192 15048
rect 22244 15036 22250 15088
rect 22094 15017 22100 15020
rect 21821 15011 21879 15017
rect 21821 14977 21833 15011
rect 21867 14977 21879 15011
rect 21821 14971 21879 14977
rect 22088 14971 22100 15017
rect 22152 15008 22158 15020
rect 23584 15008 23612 15116
rect 32858 15104 32864 15156
rect 32916 15144 32922 15156
rect 33134 15144 33140 15156
rect 32916 15116 33140 15144
rect 32916 15104 32922 15116
rect 33134 15104 33140 15116
rect 33192 15104 33198 15156
rect 33410 15104 33416 15156
rect 33468 15144 33474 15156
rect 34057 15147 34115 15153
rect 34057 15144 34069 15147
rect 33468 15116 34069 15144
rect 33468 15104 33474 15116
rect 34057 15113 34069 15116
rect 34103 15113 34115 15147
rect 36357 15147 36415 15153
rect 36357 15144 36369 15147
rect 34057 15107 34115 15113
rect 34624 15116 36369 15144
rect 30466 15036 30472 15088
rect 30524 15076 30530 15088
rect 32944 15079 33002 15085
rect 30524 15048 30880 15076
rect 30524 15036 30530 15048
rect 23661 15011 23719 15017
rect 23661 15008 23673 15011
rect 22152 14980 22188 15008
rect 23584 14980 23673 15008
rect 22094 14968 22100 14971
rect 22152 14968 22158 14980
rect 23661 14977 23673 14980
rect 23707 14977 23719 15011
rect 23842 15008 23848 15020
rect 23803 14980 23848 15008
rect 23661 14971 23719 14977
rect 19334 14900 19340 14952
rect 19392 14940 19398 14952
rect 19705 14943 19763 14949
rect 19705 14940 19717 14943
rect 19392 14912 19717 14940
rect 19392 14900 19398 14912
rect 19705 14909 19717 14912
rect 19751 14940 19763 14943
rect 20530 14940 20536 14952
rect 19751 14912 20536 14940
rect 19751 14909 19763 14912
rect 19705 14903 19763 14909
rect 20530 14900 20536 14912
rect 20588 14900 20594 14952
rect 23676 14940 23704 14971
rect 23842 14968 23848 14980
rect 23900 14968 23906 15020
rect 24029 15011 24087 15017
rect 24029 14977 24041 15011
rect 24075 15008 24087 15011
rect 24673 15011 24731 15017
rect 24673 15008 24685 15011
rect 24075 14980 24685 15008
rect 24075 14977 24087 14980
rect 24029 14971 24087 14977
rect 24673 14977 24685 14980
rect 24719 14977 24731 15011
rect 25590 15008 25596 15020
rect 25551 14980 25596 15008
rect 24673 14971 24731 14977
rect 25590 14968 25596 14980
rect 25648 14968 25654 15020
rect 26142 14968 26148 15020
rect 26200 15008 26206 15020
rect 28442 15008 28448 15020
rect 26200 14980 28448 15008
rect 26200 14968 26206 14980
rect 28442 14968 28448 14980
rect 28500 15008 28506 15020
rect 28629 15011 28687 15017
rect 28629 15008 28641 15011
rect 28500 14980 28641 15008
rect 28500 14968 28506 14980
rect 28629 14977 28641 14980
rect 28675 14977 28687 15011
rect 28629 14971 28687 14977
rect 28813 15011 28871 15017
rect 28813 14977 28825 15011
rect 28859 15008 28871 15011
rect 28994 15008 29000 15020
rect 28859 14980 29000 15008
rect 28859 14977 28871 14980
rect 28813 14971 28871 14977
rect 28994 14968 29000 14980
rect 29052 14968 29058 15020
rect 30009 15011 30067 15017
rect 30009 14977 30021 15011
rect 30055 15008 30067 15011
rect 30558 15008 30564 15020
rect 30055 14980 30564 15008
rect 30055 14977 30067 14980
rect 30009 14971 30067 14977
rect 30558 14968 30564 14980
rect 30616 14968 30622 15020
rect 30852 15017 30880 15048
rect 32944 15045 32956 15079
rect 32990 15076 33002 15079
rect 34624 15076 34652 15116
rect 36357 15113 36369 15116
rect 36403 15113 36415 15147
rect 36357 15107 36415 15113
rect 34773 15079 34831 15085
rect 34773 15076 34785 15079
rect 32990 15048 34652 15076
rect 34716 15048 34785 15076
rect 32990 15045 33002 15048
rect 32944 15039 33002 15045
rect 30837 15011 30895 15017
rect 30837 14977 30849 15011
rect 30883 14977 30895 15011
rect 34422 15008 34428 15020
rect 30837 14971 30895 14977
rect 32692 14980 34428 15008
rect 32692 14952 32720 14980
rect 34422 14968 34428 14980
rect 34480 15008 34486 15020
rect 34517 15011 34575 15017
rect 34517 15008 34529 15011
rect 34480 14980 34529 15008
rect 34480 14968 34486 14980
rect 34517 14977 34529 14980
rect 34563 14977 34575 15011
rect 34716 15008 34744 15048
rect 34773 15045 34785 15048
rect 34819 15045 34831 15079
rect 34773 15039 34831 15045
rect 34517 14971 34575 14977
rect 34624 14980 34744 15008
rect 25409 14943 25467 14949
rect 25409 14940 25421 14943
rect 23676 14912 25421 14940
rect 25409 14909 25421 14912
rect 25455 14940 25467 14943
rect 29825 14943 29883 14949
rect 29825 14940 29837 14943
rect 25455 14912 29837 14940
rect 25455 14909 25467 14912
rect 25409 14903 25467 14909
rect 29825 14909 29837 14912
rect 29871 14940 29883 14943
rect 30653 14943 30711 14949
rect 30653 14940 30665 14943
rect 29871 14912 30665 14940
rect 29871 14909 29883 14912
rect 29825 14903 29883 14909
rect 30653 14909 30665 14912
rect 30699 14909 30711 14943
rect 32674 14940 32680 14952
rect 32587 14912 32680 14940
rect 30653 14903 30711 14909
rect 32674 14900 32680 14912
rect 32732 14900 32738 14952
rect 33962 14900 33968 14952
rect 34020 14940 34026 14952
rect 34624 14940 34652 14980
rect 35802 14968 35808 15020
rect 35860 15008 35866 15020
rect 36541 15011 36599 15017
rect 36541 15008 36553 15011
rect 35860 14980 36553 15008
rect 35860 14968 35866 14980
rect 36541 14977 36553 14980
rect 36587 14977 36599 15011
rect 36541 14971 36599 14977
rect 34020 14912 34652 14940
rect 34020 14900 34026 14912
rect 29546 14832 29552 14884
rect 29604 14872 29610 14884
rect 32692 14872 32720 14900
rect 29604 14844 32720 14872
rect 33796 14844 34192 14872
rect 29604 14832 29610 14844
rect 18064 14776 19288 14804
rect 19426 14764 19432 14816
rect 19484 14804 19490 14816
rect 20162 14804 20168 14816
rect 19484 14776 20168 14804
rect 19484 14764 19490 14776
rect 20162 14764 20168 14776
rect 20220 14764 20226 14816
rect 22002 14764 22008 14816
rect 22060 14804 22066 14816
rect 23201 14807 23259 14813
rect 23201 14804 23213 14807
rect 22060 14776 23213 14804
rect 22060 14764 22066 14776
rect 23201 14773 23213 14776
rect 23247 14773 23259 14807
rect 23201 14767 23259 14773
rect 24302 14764 24308 14816
rect 24360 14804 24366 14816
rect 24489 14807 24547 14813
rect 24489 14804 24501 14807
rect 24360 14776 24501 14804
rect 24360 14764 24366 14776
rect 24489 14773 24501 14776
rect 24535 14773 24547 14807
rect 24489 14767 24547 14773
rect 25777 14807 25835 14813
rect 25777 14773 25789 14807
rect 25823 14804 25835 14807
rect 26602 14804 26608 14816
rect 25823 14776 26608 14804
rect 25823 14773 25835 14776
rect 25777 14767 25835 14773
rect 26602 14764 26608 14776
rect 26660 14764 26666 14816
rect 28629 14807 28687 14813
rect 28629 14773 28641 14807
rect 28675 14804 28687 14807
rect 29638 14804 29644 14816
rect 28675 14776 29644 14804
rect 28675 14773 28687 14776
rect 28629 14767 28687 14773
rect 29638 14764 29644 14776
rect 29696 14764 29702 14816
rect 29914 14764 29920 14816
rect 29972 14804 29978 14816
rect 30193 14807 30251 14813
rect 30193 14804 30205 14807
rect 29972 14776 30205 14804
rect 29972 14764 29978 14776
rect 30193 14773 30205 14776
rect 30239 14773 30251 14807
rect 30193 14767 30251 14773
rect 31021 14807 31079 14813
rect 31021 14773 31033 14807
rect 31067 14804 31079 14807
rect 31570 14804 31576 14816
rect 31067 14776 31576 14804
rect 31067 14773 31079 14776
rect 31021 14767 31079 14773
rect 31570 14764 31576 14776
rect 31628 14764 31634 14816
rect 31846 14764 31852 14816
rect 31904 14804 31910 14816
rect 33796 14804 33824 14844
rect 31904 14776 33824 14804
rect 34164 14804 34192 14844
rect 35897 14807 35955 14813
rect 35897 14804 35909 14807
rect 34164 14776 35909 14804
rect 31904 14764 31910 14776
rect 35897 14773 35909 14776
rect 35943 14773 35955 14807
rect 35897 14767 35955 14773
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 3237 14603 3295 14609
rect 3237 14569 3249 14603
rect 3283 14600 3295 14603
rect 4706 14600 4712 14612
rect 3283 14572 4712 14600
rect 3283 14569 3295 14572
rect 3237 14563 3295 14569
rect 4706 14560 4712 14572
rect 4764 14560 4770 14612
rect 8110 14560 8116 14612
rect 8168 14600 8174 14612
rect 8205 14603 8263 14609
rect 8205 14600 8217 14603
rect 8168 14572 8217 14600
rect 8168 14560 8174 14572
rect 8205 14569 8217 14572
rect 8251 14569 8263 14603
rect 8205 14563 8263 14569
rect 12434 14560 12440 14612
rect 12492 14600 12498 14612
rect 13449 14603 13507 14609
rect 13449 14600 13461 14603
rect 12492 14572 13461 14600
rect 12492 14560 12498 14572
rect 13449 14569 13461 14572
rect 13495 14600 13507 14603
rect 14826 14600 14832 14612
rect 13495 14572 14832 14600
rect 13495 14569 13507 14572
rect 13449 14563 13507 14569
rect 14826 14560 14832 14572
rect 14884 14560 14890 14612
rect 18322 14560 18328 14612
rect 18380 14600 18386 14612
rect 20070 14600 20076 14612
rect 18380 14572 20076 14600
rect 18380 14560 18386 14572
rect 20070 14560 20076 14572
rect 20128 14560 20134 14612
rect 20438 14560 20444 14612
rect 20496 14600 20502 14612
rect 20898 14600 20904 14612
rect 20496 14572 20904 14600
rect 20496 14560 20502 14572
rect 20898 14560 20904 14572
rect 20956 14560 20962 14612
rect 21910 14560 21916 14612
rect 21968 14600 21974 14612
rect 22005 14603 22063 14609
rect 22005 14600 22017 14603
rect 21968 14572 22017 14600
rect 21968 14560 21974 14572
rect 22005 14569 22017 14572
rect 22051 14569 22063 14603
rect 22005 14563 22063 14569
rect 24854 14560 24860 14612
rect 24912 14600 24918 14612
rect 26053 14603 26111 14609
rect 26053 14600 26065 14603
rect 24912 14572 26065 14600
rect 24912 14560 24918 14572
rect 26053 14569 26065 14572
rect 26099 14569 26111 14603
rect 26053 14563 26111 14569
rect 27890 14560 27896 14612
rect 27948 14600 27954 14612
rect 28077 14603 28135 14609
rect 28077 14600 28089 14603
rect 27948 14572 28089 14600
rect 27948 14560 27954 14572
rect 28077 14569 28089 14572
rect 28123 14600 28135 14603
rect 28813 14603 28871 14609
rect 28813 14600 28825 14603
rect 28123 14572 28825 14600
rect 28123 14569 28135 14572
rect 28077 14563 28135 14569
rect 28813 14569 28825 14572
rect 28859 14569 28871 14603
rect 28994 14600 29000 14612
rect 28813 14563 28871 14569
rect 28920 14572 29000 14600
rect 5350 14492 5356 14544
rect 5408 14532 5414 14544
rect 15562 14532 15568 14544
rect 5408 14504 8248 14532
rect 5408 14492 5414 14504
rect 8220 14476 8248 14504
rect 13832 14504 15568 14532
rect 3786 14464 3792 14476
rect 3747 14436 3792 14464
rect 3786 14424 3792 14436
rect 3844 14424 3850 14476
rect 6178 14464 6184 14476
rect 4816 14436 6184 14464
rect 1857 14399 1915 14405
rect 1857 14365 1869 14399
rect 1903 14396 1915 14399
rect 2682 14396 2688 14408
rect 1903 14368 2688 14396
rect 1903 14365 1915 14368
rect 1857 14359 1915 14365
rect 2682 14356 2688 14368
rect 2740 14396 2746 14408
rect 3804 14396 3832 14424
rect 2740 14368 3832 14396
rect 4056 14399 4114 14405
rect 2740 14356 2746 14368
rect 4056 14365 4068 14399
rect 4102 14396 4114 14399
rect 4614 14396 4620 14408
rect 4102 14368 4620 14396
rect 4102 14365 4114 14368
rect 4056 14359 4114 14365
rect 4614 14356 4620 14368
rect 4672 14356 4678 14408
rect 2124 14331 2182 14337
rect 2124 14297 2136 14331
rect 2170 14328 2182 14331
rect 4816 14328 4844 14436
rect 6178 14424 6184 14436
rect 6236 14424 6242 14476
rect 8202 14424 8208 14476
rect 8260 14424 8266 14476
rect 9766 14464 9772 14476
rect 9727 14436 9772 14464
rect 9766 14424 9772 14436
rect 9824 14424 9830 14476
rect 5629 14399 5687 14405
rect 5629 14365 5641 14399
rect 5675 14396 5687 14399
rect 8386 14396 8392 14408
rect 5675 14368 8392 14396
rect 5675 14365 5687 14368
rect 5629 14359 5687 14365
rect 8386 14356 8392 14368
rect 8444 14356 8450 14408
rect 9122 14396 9128 14408
rect 9083 14368 9128 14396
rect 9122 14356 9128 14368
rect 9180 14356 9186 14408
rect 12066 14396 12072 14408
rect 12027 14368 12072 14396
rect 12066 14356 12072 14368
rect 12124 14356 12130 14408
rect 2170 14300 4844 14328
rect 5184 14300 7788 14328
rect 2170 14297 2182 14300
rect 2124 14291 2182 14297
rect 5184 14269 5212 14300
rect 5169 14263 5227 14269
rect 5169 14229 5181 14263
rect 5215 14229 5227 14263
rect 5169 14223 5227 14229
rect 6822 14220 6828 14272
rect 6880 14260 6886 14272
rect 6917 14263 6975 14269
rect 6917 14260 6929 14263
rect 6880 14232 6929 14260
rect 6880 14220 6886 14232
rect 6917 14229 6929 14232
rect 6963 14229 6975 14263
rect 7760 14260 7788 14300
rect 7834 14288 7840 14340
rect 7892 14328 7898 14340
rect 8021 14331 8079 14337
rect 7892 14300 7937 14328
rect 7892 14288 7898 14300
rect 8021 14297 8033 14331
rect 8067 14297 8079 14331
rect 8021 14291 8079 14297
rect 10036 14331 10094 14337
rect 10036 14297 10048 14331
rect 10082 14328 10094 14331
rect 11606 14328 11612 14340
rect 10082 14300 11612 14328
rect 10082 14297 10094 14300
rect 10036 14291 10094 14297
rect 8036 14260 8064 14291
rect 11606 14288 11612 14300
rect 11664 14288 11670 14340
rect 12336 14331 12394 14337
rect 12336 14297 12348 14331
rect 12382 14328 12394 14331
rect 13170 14328 13176 14340
rect 12382 14300 13176 14328
rect 12382 14297 12394 14300
rect 12336 14291 12394 14297
rect 13170 14288 13176 14300
rect 13228 14288 13234 14340
rect 8938 14260 8944 14272
rect 7760 14232 8064 14260
rect 8899 14232 8944 14260
rect 6917 14223 6975 14229
rect 8938 14220 8944 14232
rect 8996 14220 9002 14272
rect 10318 14220 10324 14272
rect 10376 14260 10382 14272
rect 11149 14263 11207 14269
rect 11149 14260 11161 14263
rect 10376 14232 11161 14260
rect 10376 14220 10382 14232
rect 11149 14229 11161 14232
rect 11195 14260 11207 14263
rect 13832 14260 13860 14504
rect 15562 14492 15568 14504
rect 15620 14492 15626 14544
rect 16301 14535 16359 14541
rect 16301 14501 16313 14535
rect 16347 14532 16359 14535
rect 16482 14532 16488 14544
rect 16347 14504 16488 14532
rect 16347 14501 16359 14504
rect 16301 14495 16359 14501
rect 16482 14492 16488 14504
rect 16540 14492 16546 14544
rect 23014 14532 23020 14544
rect 19168 14504 23020 14532
rect 15194 14424 15200 14476
rect 15252 14464 15258 14476
rect 15252 14436 15792 14464
rect 15252 14424 15258 14436
rect 15105 14399 15163 14405
rect 15105 14365 15117 14399
rect 15151 14365 15163 14399
rect 15378 14396 15384 14408
rect 15339 14368 15384 14396
rect 15105 14359 15163 14365
rect 15120 14328 15148 14359
rect 15378 14356 15384 14368
rect 15436 14356 15442 14408
rect 15764 14405 15792 14436
rect 16206 14424 16212 14476
rect 16264 14464 16270 14476
rect 16264 14436 18184 14464
rect 16264 14424 16270 14436
rect 15749 14399 15807 14405
rect 15749 14365 15761 14399
rect 15795 14365 15807 14399
rect 15749 14359 15807 14365
rect 16301 14399 16359 14405
rect 16301 14365 16313 14399
rect 16347 14396 16359 14399
rect 16666 14396 16672 14408
rect 16347 14368 16672 14396
rect 16347 14365 16359 14368
rect 16301 14359 16359 14365
rect 16666 14356 16672 14368
rect 16724 14356 16730 14408
rect 17494 14396 17500 14408
rect 17455 14368 17500 14396
rect 17494 14356 17500 14368
rect 17552 14356 17558 14408
rect 17862 14396 17868 14408
rect 17823 14368 17868 14396
rect 17862 14356 17868 14368
rect 17920 14356 17926 14408
rect 18049 14399 18107 14405
rect 18049 14365 18061 14399
rect 18095 14365 18107 14399
rect 18049 14359 18107 14365
rect 15654 14328 15660 14340
rect 15120 14300 15660 14328
rect 15654 14288 15660 14300
rect 15712 14288 15718 14340
rect 16850 14288 16856 14340
rect 16908 14328 16914 14340
rect 18064 14328 18092 14359
rect 16908 14300 18092 14328
rect 18156 14328 18184 14436
rect 18325 14399 18383 14405
rect 18325 14365 18337 14399
rect 18371 14396 18383 14399
rect 19168 14396 19196 14504
rect 23014 14492 23020 14504
rect 23072 14492 23078 14544
rect 28920 14541 28948 14572
rect 28994 14560 29000 14572
rect 29052 14560 29058 14612
rect 33781 14603 33839 14609
rect 33781 14569 33793 14603
rect 33827 14600 33839 14603
rect 34606 14600 34612 14612
rect 33827 14572 34612 14600
rect 33827 14569 33839 14572
rect 33781 14563 33839 14569
rect 34606 14560 34612 14572
rect 34664 14560 34670 14612
rect 35894 14600 35900 14612
rect 34716 14572 35900 14600
rect 28905 14535 28963 14541
rect 28905 14501 28917 14535
rect 28951 14501 28963 14535
rect 34716 14532 34744 14572
rect 35894 14560 35900 14572
rect 35952 14560 35958 14612
rect 28905 14495 28963 14501
rect 32324 14504 34744 14532
rect 26142 14464 26148 14476
rect 19260 14436 26148 14464
rect 19260 14405 19288 14436
rect 26142 14424 26148 14436
rect 26200 14424 26206 14476
rect 28258 14464 28264 14476
rect 28219 14436 28264 14464
rect 28258 14424 28264 14436
rect 28316 14424 28322 14476
rect 18371 14368 19196 14396
rect 19245 14399 19303 14405
rect 18371 14365 18383 14368
rect 18325 14359 18383 14365
rect 19245 14365 19257 14399
rect 19291 14365 19303 14399
rect 19245 14359 19303 14365
rect 19260 14328 19288 14359
rect 19334 14356 19340 14408
rect 19392 14396 19398 14408
rect 19521 14399 19579 14405
rect 19521 14396 19533 14399
rect 19392 14368 19533 14396
rect 19392 14356 19398 14368
rect 19521 14365 19533 14368
rect 19567 14365 19579 14399
rect 19521 14359 19579 14365
rect 19981 14399 20039 14405
rect 19981 14365 19993 14399
rect 20027 14396 20039 14399
rect 20070 14396 20076 14408
rect 20027 14368 20076 14396
rect 20027 14365 20039 14368
rect 19981 14359 20039 14365
rect 19426 14328 19432 14340
rect 18156 14300 19288 14328
rect 19339 14300 19432 14328
rect 16908 14288 16914 14300
rect 19426 14288 19432 14300
rect 19484 14328 19490 14340
rect 19996 14328 20024 14359
rect 20070 14356 20076 14368
rect 20128 14356 20134 14408
rect 20165 14399 20223 14405
rect 20165 14365 20177 14399
rect 20211 14396 20223 14399
rect 20438 14396 20444 14408
rect 20211 14368 20444 14396
rect 20211 14365 20223 14368
rect 20165 14359 20223 14365
rect 20438 14356 20444 14368
rect 20496 14356 20502 14408
rect 21913 14399 21971 14405
rect 21913 14365 21925 14399
rect 21959 14396 21971 14399
rect 22002 14396 22008 14408
rect 21959 14368 22008 14396
rect 21959 14365 21971 14368
rect 21913 14359 21971 14365
rect 22002 14356 22008 14368
rect 22060 14356 22066 14408
rect 22738 14356 22744 14408
rect 22796 14396 22802 14408
rect 23201 14399 23259 14405
rect 23201 14396 23213 14399
rect 22796 14368 23213 14396
rect 22796 14356 22802 14368
rect 23201 14365 23213 14368
rect 23247 14365 23259 14399
rect 26970 14396 26976 14408
rect 26931 14368 26976 14396
rect 23201 14359 23259 14365
rect 26970 14356 26976 14368
rect 27028 14356 27034 14408
rect 27154 14396 27160 14408
rect 27115 14368 27160 14396
rect 27154 14356 27160 14368
rect 27212 14356 27218 14408
rect 27982 14396 27988 14408
rect 27943 14368 27988 14396
rect 27982 14356 27988 14368
rect 28040 14356 28046 14408
rect 28721 14399 28779 14405
rect 28721 14365 28733 14399
rect 28767 14365 28779 14399
rect 28920 14396 28948 14495
rect 28997 14467 29055 14473
rect 28997 14433 29009 14467
rect 29043 14464 29055 14467
rect 29086 14464 29092 14476
rect 29043 14436 29092 14464
rect 29043 14433 29055 14436
rect 28997 14427 29055 14433
rect 29086 14424 29092 14436
rect 29144 14424 29150 14476
rect 29546 14464 29552 14476
rect 29507 14436 29552 14464
rect 29546 14424 29552 14436
rect 29604 14424 29610 14476
rect 28920 14368 29592 14396
rect 28721 14359 28779 14365
rect 23934 14328 23940 14340
rect 19484 14300 19564 14328
rect 19996 14300 23940 14328
rect 19484 14288 19490 14300
rect 11195 14232 13860 14260
rect 11195 14229 11207 14232
rect 11149 14223 11207 14229
rect 15102 14220 15108 14272
rect 15160 14260 15166 14272
rect 17402 14260 17408 14272
rect 15160 14232 17408 14260
rect 15160 14220 15166 14232
rect 17402 14220 17408 14232
rect 17460 14220 17466 14272
rect 19334 14260 19340 14272
rect 19392 14269 19398 14272
rect 19301 14232 19340 14260
rect 19334 14220 19340 14232
rect 19392 14223 19401 14269
rect 19536 14260 19564 14300
rect 23934 14288 23940 14300
rect 23992 14288 23998 14340
rect 24762 14328 24768 14340
rect 24723 14300 24768 14328
rect 24762 14288 24768 14300
rect 24820 14288 24826 14340
rect 26988 14328 27016 14356
rect 27522 14328 27528 14340
rect 26988 14300 27528 14328
rect 27522 14288 27528 14300
rect 27580 14288 27586 14340
rect 28736 14328 28764 14359
rect 29564 14340 29592 14368
rect 29638 14356 29644 14408
rect 29696 14396 29702 14408
rect 29805 14399 29863 14405
rect 29805 14396 29817 14399
rect 29696 14368 29817 14396
rect 29696 14356 29702 14368
rect 29805 14365 29817 14368
rect 29851 14365 29863 14399
rect 31570 14396 31576 14408
rect 31531 14368 31576 14396
rect 29805 14359 29863 14365
rect 31570 14356 31576 14368
rect 31628 14356 31634 14408
rect 32324 14405 32352 14504
rect 32674 14424 32680 14476
rect 32732 14464 32738 14476
rect 32732 14436 34100 14464
rect 32732 14424 32738 14436
rect 32309 14399 32367 14405
rect 32309 14365 32321 14399
rect 32355 14365 32367 14399
rect 32309 14359 32367 14365
rect 32493 14399 32551 14405
rect 32493 14365 32505 14399
rect 32539 14396 32551 14399
rect 33965 14399 34023 14405
rect 33965 14396 33977 14399
rect 32539 14368 33977 14396
rect 32539 14365 32551 14368
rect 32493 14359 32551 14365
rect 33965 14365 33977 14368
rect 34011 14365 34023 14399
rect 34072 14396 34100 14436
rect 34422 14424 34428 14476
rect 34480 14464 34486 14476
rect 34701 14467 34759 14473
rect 34701 14464 34713 14467
rect 34480 14436 34713 14464
rect 34480 14424 34486 14436
rect 34701 14433 34713 14436
rect 34747 14433 34759 14467
rect 34701 14427 34759 14433
rect 34072 14368 34652 14396
rect 33965 14359 34023 14365
rect 28736 14300 29132 14328
rect 20073 14263 20131 14269
rect 20073 14260 20085 14263
rect 19536 14232 20085 14260
rect 20073 14229 20085 14232
rect 20119 14229 20131 14263
rect 20073 14223 20131 14229
rect 19392 14220 19398 14223
rect 20898 14220 20904 14272
rect 20956 14260 20962 14272
rect 23106 14260 23112 14272
rect 20956 14232 23112 14260
rect 20956 14220 20962 14232
rect 23106 14220 23112 14232
rect 23164 14260 23170 14272
rect 23385 14263 23443 14269
rect 23385 14260 23397 14263
rect 23164 14232 23397 14260
rect 23164 14220 23170 14232
rect 23385 14229 23397 14232
rect 23431 14229 23443 14263
rect 27062 14260 27068 14272
rect 27023 14232 27068 14260
rect 23385 14223 23443 14229
rect 27062 14220 27068 14232
rect 27120 14220 27126 14272
rect 28258 14260 28264 14272
rect 28219 14232 28264 14260
rect 28258 14220 28264 14232
rect 28316 14220 28322 14272
rect 29104 14260 29132 14300
rect 29546 14288 29552 14340
rect 29604 14288 29610 14340
rect 32122 14328 32128 14340
rect 32083 14300 32128 14328
rect 32122 14288 32128 14300
rect 32180 14288 32186 14340
rect 32398 14288 32404 14340
rect 32456 14328 32462 14340
rect 32766 14328 32772 14340
rect 32456 14300 32772 14328
rect 32456 14288 32462 14300
rect 32766 14288 32772 14300
rect 32824 14328 32830 14340
rect 32953 14331 33011 14337
rect 32953 14328 32965 14331
rect 32824 14300 32965 14328
rect 32824 14288 32830 14300
rect 32953 14297 32965 14300
rect 32999 14297 33011 14331
rect 32953 14291 33011 14297
rect 33137 14331 33195 14337
rect 33137 14297 33149 14331
rect 33183 14328 33195 14331
rect 34514 14328 34520 14340
rect 33183 14300 34520 14328
rect 33183 14297 33195 14300
rect 33137 14291 33195 14297
rect 34514 14288 34520 14300
rect 34572 14288 34578 14340
rect 34624 14328 34652 14368
rect 34790 14356 34796 14408
rect 34848 14396 34854 14408
rect 34957 14399 35015 14405
rect 34957 14396 34969 14399
rect 34848 14368 34969 14396
rect 34848 14356 34854 14368
rect 34957 14365 34969 14368
rect 35003 14365 35015 14399
rect 34957 14359 35015 14365
rect 36078 14356 36084 14408
rect 36136 14356 36142 14408
rect 36096 14328 36124 14356
rect 34624 14300 36124 14328
rect 30929 14263 30987 14269
rect 30929 14260 30941 14263
rect 29104 14232 30941 14260
rect 30929 14229 30941 14232
rect 30975 14229 30987 14263
rect 30929 14223 30987 14229
rect 31389 14263 31447 14269
rect 31389 14229 31401 14263
rect 31435 14260 31447 14263
rect 32030 14260 32036 14272
rect 31435 14232 32036 14260
rect 31435 14229 31447 14232
rect 31389 14223 31447 14229
rect 32030 14220 32036 14232
rect 32088 14220 32094 14272
rect 33318 14260 33324 14272
rect 33279 14232 33324 14260
rect 33318 14220 33324 14232
rect 33376 14220 33382 14272
rect 33410 14220 33416 14272
rect 33468 14260 33474 14272
rect 36081 14263 36139 14269
rect 36081 14260 36093 14263
rect 33468 14232 36093 14260
rect 33468 14220 33474 14232
rect 36081 14229 36093 14232
rect 36127 14229 36139 14263
rect 36081 14223 36139 14229
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 4065 14059 4123 14065
rect 4065 14025 4077 14059
rect 4111 14056 4123 14059
rect 5626 14056 5632 14068
rect 4111 14028 5632 14056
rect 4111 14025 4123 14028
rect 4065 14019 4123 14025
rect 5626 14016 5632 14028
rect 5684 14016 5690 14068
rect 6270 14016 6276 14068
rect 6328 14056 6334 14068
rect 6733 14059 6791 14065
rect 6733 14056 6745 14059
rect 6328 14028 6745 14056
rect 6328 14016 6334 14028
rect 6733 14025 6745 14028
rect 6779 14025 6791 14059
rect 6733 14019 6791 14025
rect 7098 14016 7104 14068
rect 7156 14056 7162 14068
rect 7561 14059 7619 14065
rect 7561 14056 7573 14059
rect 7156 14028 7573 14056
rect 7156 14016 7162 14028
rect 7561 14025 7573 14028
rect 7607 14025 7619 14059
rect 11606 14056 11612 14068
rect 11567 14028 11612 14056
rect 7561 14019 7619 14025
rect 11606 14016 11612 14028
rect 11664 14016 11670 14068
rect 13170 14056 13176 14068
rect 13131 14028 13176 14056
rect 13170 14016 13176 14028
rect 13228 14016 13234 14068
rect 14185 14059 14243 14065
rect 14185 14025 14197 14059
rect 14231 14056 14243 14059
rect 15378 14056 15384 14068
rect 14231 14028 15384 14056
rect 14231 14025 14243 14028
rect 14185 14019 14243 14025
rect 15378 14016 15384 14028
rect 15436 14016 15442 14068
rect 16025 14059 16083 14065
rect 16025 14025 16037 14059
rect 16071 14056 16083 14059
rect 18046 14056 18052 14068
rect 16071 14028 18052 14056
rect 16071 14025 16083 14028
rect 16025 14019 16083 14025
rect 18046 14016 18052 14028
rect 18104 14016 18110 14068
rect 20438 14056 20444 14068
rect 20399 14028 20444 14056
rect 20438 14016 20444 14028
rect 20496 14016 20502 14068
rect 24762 14016 24768 14068
rect 24820 14056 24826 14068
rect 29733 14059 29791 14065
rect 24820 14028 28994 14056
rect 24820 14016 24826 14028
rect 2952 13991 3010 13997
rect 2952 13957 2964 13991
rect 2998 13988 3010 13991
rect 4798 13988 4804 14000
rect 2998 13960 4804 13988
rect 2998 13957 3010 13960
rect 2952 13951 3010 13957
rect 4798 13948 4804 13960
rect 4856 13948 4862 14000
rect 6638 13988 6644 14000
rect 5828 13960 6644 13988
rect 2682 13920 2688 13932
rect 2643 13892 2688 13920
rect 2682 13880 2688 13892
rect 2740 13880 2746 13932
rect 5828 13929 5856 13960
rect 6638 13948 6644 13960
rect 6696 13948 6702 14000
rect 7006 13948 7012 14000
rect 7064 13988 7070 14000
rect 7377 13991 7435 13997
rect 7377 13988 7389 13991
rect 7064 13960 7389 13988
rect 7064 13948 7070 13960
rect 7377 13957 7389 13960
rect 7423 13957 7435 13991
rect 7377 13951 7435 13957
rect 8110 13948 8116 14000
rect 8168 13988 8174 14000
rect 9401 13991 9459 13997
rect 9401 13988 9413 13991
rect 8168 13960 9413 13988
rect 8168 13948 8174 13960
rect 9401 13957 9413 13960
rect 9447 13957 9459 13991
rect 9401 13951 9459 13957
rect 10042 13948 10048 14000
rect 10100 13988 10106 14000
rect 10137 13991 10195 13997
rect 10137 13988 10149 13991
rect 10100 13960 10149 13988
rect 10100 13948 10106 13960
rect 10137 13957 10149 13960
rect 10183 13988 10195 13991
rect 12158 13988 12164 14000
rect 10183 13960 12164 13988
rect 10183 13957 10195 13960
rect 10137 13951 10195 13957
rect 12158 13948 12164 13960
rect 12216 13948 12222 14000
rect 12323 13991 12381 13997
rect 12323 13957 12335 13991
rect 12369 13988 12381 13991
rect 15654 13988 15660 14000
rect 12369 13960 13032 13988
rect 12369 13957 12381 13960
rect 12323 13951 12381 13957
rect 5813 13923 5871 13929
rect 5813 13889 5825 13923
rect 5859 13889 5871 13923
rect 6362 13920 6368 13932
rect 6275 13892 6368 13920
rect 5813 13883 5871 13889
rect 6362 13880 6368 13892
rect 6420 13880 6426 13932
rect 6546 13920 6552 13932
rect 6507 13892 6552 13920
rect 6546 13880 6552 13892
rect 6604 13880 6610 13932
rect 7190 13920 7196 13932
rect 7151 13892 7196 13920
rect 7190 13880 7196 13892
rect 7248 13920 7254 13932
rect 7834 13920 7840 13932
rect 7248 13892 7840 13920
rect 7248 13880 7254 13892
rect 7834 13880 7840 13892
rect 7892 13880 7898 13932
rect 8202 13920 8208 13932
rect 8163 13892 8208 13920
rect 8202 13880 8208 13892
rect 8260 13880 8266 13932
rect 8294 13880 8300 13932
rect 8352 13920 8358 13932
rect 8389 13923 8447 13929
rect 8389 13920 8401 13923
rect 8352 13892 8401 13920
rect 8352 13880 8358 13892
rect 8389 13889 8401 13892
rect 8435 13889 8447 13923
rect 9033 13923 9091 13929
rect 9033 13920 9045 13923
rect 8389 13883 8447 13889
rect 8496 13892 9045 13920
rect 5718 13852 5724 13864
rect 5644 13824 5724 13852
rect 5644 13793 5672 13824
rect 5718 13812 5724 13824
rect 5776 13812 5782 13864
rect 6380 13852 6408 13880
rect 6730 13852 6736 13864
rect 6380 13824 6736 13852
rect 6730 13812 6736 13824
rect 6788 13812 6794 13864
rect 7852 13852 7880 13880
rect 8496 13852 8524 13892
rect 9033 13889 9045 13892
rect 9079 13889 9091 13923
rect 9214 13920 9220 13932
rect 9175 13892 9220 13920
rect 9033 13883 9091 13889
rect 9214 13880 9220 13892
rect 9272 13880 9278 13932
rect 10502 13920 10508 13932
rect 10463 13892 10508 13920
rect 10502 13880 10508 13892
rect 10560 13880 10566 13932
rect 11517 13923 11575 13929
rect 11517 13920 11529 13923
rect 10980 13892 11529 13920
rect 7852 13824 8524 13852
rect 8573 13855 8631 13861
rect 8573 13821 8585 13855
rect 8619 13852 8631 13855
rect 9766 13852 9772 13864
rect 8619 13824 9772 13852
rect 8619 13821 8631 13824
rect 8573 13815 8631 13821
rect 9766 13812 9772 13824
rect 9824 13812 9830 13864
rect 10318 13852 10324 13864
rect 10279 13824 10324 13852
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 5629 13787 5687 13793
rect 5629 13753 5641 13787
rect 5675 13753 5687 13787
rect 10980 13784 11008 13892
rect 11517 13889 11529 13892
rect 11563 13889 11575 13923
rect 11517 13883 11575 13889
rect 11701 13923 11759 13929
rect 11701 13889 11713 13923
rect 11747 13920 11759 13923
rect 11790 13920 11796 13932
rect 11747 13892 11796 13920
rect 11747 13889 11759 13892
rect 11701 13883 11759 13889
rect 11790 13880 11796 13892
rect 11848 13880 11854 13932
rect 12621 13923 12679 13929
rect 12621 13889 12633 13923
rect 12667 13889 12679 13923
rect 13004 13920 13032 13960
rect 14936 13960 15660 13988
rect 13081 13923 13139 13929
rect 13081 13920 13093 13923
rect 13004 13892 13093 13920
rect 12621 13883 12679 13889
rect 13081 13889 13093 13892
rect 13127 13889 13139 13923
rect 13262 13920 13268 13932
rect 13223 13892 13268 13920
rect 13081 13883 13139 13889
rect 12434 13812 12440 13864
rect 12492 13852 12498 13864
rect 12492 13824 12537 13852
rect 12492 13812 12498 13824
rect 5629 13747 5687 13753
rect 10336 13756 11008 13784
rect 10336 13725 10364 13756
rect 12158 13744 12164 13796
rect 12216 13784 12222 13796
rect 12253 13787 12311 13793
rect 12253 13784 12265 13787
rect 12216 13756 12265 13784
rect 12216 13744 12222 13756
rect 12253 13753 12265 13756
rect 12299 13753 12311 13787
rect 12636 13784 12664 13883
rect 13262 13880 13268 13892
rect 13320 13880 13326 13932
rect 14936 13929 14964 13960
rect 15654 13948 15660 13960
rect 15712 13948 15718 14000
rect 17310 13948 17316 14000
rect 17368 13988 17374 14000
rect 19334 13997 19340 14000
rect 19328 13988 19340 13997
rect 17368 13960 19104 13988
rect 19295 13960 19340 13988
rect 17368 13948 17374 13960
rect 13817 13923 13875 13929
rect 13817 13889 13829 13923
rect 13863 13920 13875 13923
rect 14921 13923 14979 13929
rect 13863 13892 14596 13920
rect 13863 13889 13875 13892
rect 13817 13883 13875 13889
rect 13909 13855 13967 13861
rect 13909 13821 13921 13855
rect 13955 13821 13967 13855
rect 14568 13852 14596 13892
rect 14921 13889 14933 13923
rect 14967 13889 14979 13923
rect 15102 13920 15108 13932
rect 15063 13892 15108 13920
rect 14921 13883 14979 13889
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 15470 13920 15476 13932
rect 15431 13892 15476 13920
rect 15470 13880 15476 13892
rect 15528 13880 15534 13932
rect 15838 13920 15844 13932
rect 15799 13892 15844 13920
rect 15838 13880 15844 13892
rect 15896 13880 15902 13932
rect 17129 13923 17187 13929
rect 17129 13889 17141 13923
rect 17175 13889 17187 13923
rect 17129 13883 17187 13889
rect 15562 13852 15568 13864
rect 14568 13824 15568 13852
rect 13909 13815 13967 13821
rect 13170 13784 13176 13796
rect 12636 13756 13176 13784
rect 12253 13747 12311 13753
rect 13170 13744 13176 13756
rect 13228 13744 13234 13796
rect 13924 13784 13952 13815
rect 15562 13812 15568 13824
rect 15620 13812 15626 13864
rect 17144 13852 17172 13883
rect 17218 13880 17224 13932
rect 17276 13920 17282 13932
rect 19076 13929 19104 13960
rect 19328 13951 19340 13960
rect 19334 13948 19340 13951
rect 19392 13948 19398 14000
rect 22738 13988 22744 14000
rect 22112 13960 22744 13988
rect 17957 13923 18015 13929
rect 17957 13920 17969 13923
rect 17276 13892 17969 13920
rect 17276 13880 17282 13892
rect 17957 13889 17969 13892
rect 18003 13889 18015 13923
rect 17957 13883 18015 13889
rect 19061 13923 19119 13929
rect 19061 13889 19073 13923
rect 19107 13889 19119 13923
rect 19061 13883 19119 13889
rect 21542 13880 21548 13932
rect 21600 13920 21606 13932
rect 22112 13929 22140 13960
rect 22738 13948 22744 13960
rect 22796 13948 22802 14000
rect 24854 13988 24860 14000
rect 22848 13960 24860 13988
rect 21913 13923 21971 13929
rect 21913 13920 21925 13923
rect 21600 13892 21925 13920
rect 21600 13880 21606 13892
rect 21913 13889 21925 13892
rect 21959 13889 21971 13923
rect 21913 13883 21971 13889
rect 22097 13923 22155 13929
rect 22097 13889 22109 13923
rect 22143 13889 22155 13923
rect 22097 13883 22155 13889
rect 22186 13880 22192 13932
rect 22244 13920 22250 13932
rect 22848 13929 22876 13960
rect 22833 13923 22891 13929
rect 22833 13920 22845 13923
rect 22244 13892 22845 13920
rect 22244 13880 22250 13892
rect 22833 13889 22845 13892
rect 22879 13889 22891 13923
rect 22833 13883 22891 13889
rect 23100 13923 23158 13929
rect 23100 13889 23112 13923
rect 23146 13920 23158 13923
rect 23658 13920 23664 13932
rect 23146 13892 23664 13920
rect 23146 13889 23158 13892
rect 23100 13883 23158 13889
rect 23658 13880 23664 13892
rect 23716 13880 23722 13932
rect 24780 13929 24808 13960
rect 24854 13948 24860 13960
rect 24912 13988 24918 14000
rect 25590 13988 25596 14000
rect 24912 13960 25596 13988
rect 24912 13948 24918 13960
rect 25590 13948 25596 13960
rect 25648 13988 25654 14000
rect 25648 13960 27200 13988
rect 25648 13948 25654 13960
rect 24765 13923 24823 13929
rect 24765 13889 24777 13923
rect 24811 13889 24823 13923
rect 24765 13883 24823 13889
rect 25032 13923 25090 13929
rect 25032 13889 25044 13923
rect 25078 13920 25090 13923
rect 27062 13920 27068 13932
rect 25078 13892 27068 13920
rect 25078 13889 25090 13892
rect 25032 13883 25090 13889
rect 27062 13880 27068 13892
rect 27120 13880 27126 13932
rect 27172 13929 27200 13960
rect 27157 13923 27215 13929
rect 27157 13889 27169 13923
rect 27203 13889 27215 13923
rect 27157 13883 27215 13889
rect 27424 13923 27482 13929
rect 27424 13889 27436 13923
rect 27470 13920 27482 13923
rect 27706 13920 27712 13932
rect 27470 13892 27712 13920
rect 27470 13889 27482 13892
rect 27424 13883 27482 13889
rect 27706 13880 27712 13892
rect 27764 13880 27770 13932
rect 27982 13880 27988 13932
rect 28040 13920 28046 13932
rect 28040 13892 28580 13920
rect 28040 13880 28046 13892
rect 17494 13852 17500 13864
rect 17144 13824 17500 13852
rect 17494 13812 17500 13824
rect 17552 13852 17558 13864
rect 17770 13852 17776 13864
rect 17552 13824 17776 13852
rect 17552 13812 17558 13824
rect 17770 13812 17776 13824
rect 17828 13812 17834 13864
rect 17862 13812 17868 13864
rect 17920 13852 17926 13864
rect 17920 13824 17965 13852
rect 17920 13812 17926 13824
rect 20162 13812 20168 13864
rect 20220 13852 20226 13864
rect 20346 13852 20352 13864
rect 20220 13824 20352 13852
rect 20220 13812 20226 13824
rect 20346 13812 20352 13824
rect 20404 13812 20410 13864
rect 15102 13784 15108 13796
rect 13924 13756 15108 13784
rect 15102 13744 15108 13756
rect 15160 13744 15166 13796
rect 17954 13784 17960 13796
rect 17915 13756 17960 13784
rect 17954 13744 17960 13756
rect 18012 13744 18018 13796
rect 28552 13793 28580 13892
rect 28537 13787 28595 13793
rect 24136 13756 24808 13784
rect 10321 13719 10379 13725
rect 10321 13685 10333 13719
rect 10367 13685 10379 13719
rect 10321 13679 10379 13685
rect 10410 13676 10416 13728
rect 10468 13716 10474 13728
rect 12529 13719 12587 13725
rect 12529 13716 12541 13719
rect 10468 13688 12541 13716
rect 10468 13676 10474 13688
rect 12529 13685 12541 13688
rect 12575 13685 12587 13719
rect 12529 13679 12587 13685
rect 14001 13719 14059 13725
rect 14001 13685 14013 13719
rect 14047 13716 14059 13719
rect 15470 13716 15476 13728
rect 14047 13688 15476 13716
rect 14047 13685 14059 13688
rect 14001 13679 14059 13685
rect 15470 13676 15476 13688
rect 15528 13676 15534 13728
rect 22005 13719 22063 13725
rect 22005 13685 22017 13719
rect 22051 13716 22063 13719
rect 24136 13716 24164 13756
rect 22051 13688 24164 13716
rect 24213 13719 24271 13725
rect 22051 13685 22063 13688
rect 22005 13679 22063 13685
rect 24213 13685 24225 13719
rect 24259 13716 24271 13719
rect 24394 13716 24400 13728
rect 24259 13688 24400 13716
rect 24259 13685 24271 13688
rect 24213 13679 24271 13685
rect 24394 13676 24400 13688
rect 24452 13676 24458 13728
rect 24780 13716 24808 13756
rect 28537 13753 28549 13787
rect 28583 13753 28595 13787
rect 28537 13747 28595 13753
rect 26050 13716 26056 13728
rect 24780 13688 26056 13716
rect 26050 13676 26056 13688
rect 26108 13676 26114 13728
rect 26145 13719 26203 13725
rect 26145 13685 26157 13719
rect 26191 13716 26203 13719
rect 26234 13716 26240 13728
rect 26191 13688 26240 13716
rect 26191 13685 26203 13688
rect 26145 13679 26203 13685
rect 26234 13676 26240 13688
rect 26292 13676 26298 13728
rect 28966 13716 28994 14028
rect 29733 14025 29745 14059
rect 29779 14056 29791 14059
rect 30650 14056 30656 14068
rect 29779 14028 30656 14056
rect 29779 14025 29791 14028
rect 29733 14019 29791 14025
rect 30650 14016 30656 14028
rect 30708 14016 30714 14068
rect 31389 14059 31447 14065
rect 31389 14025 31401 14059
rect 31435 14056 31447 14059
rect 32858 14056 32864 14068
rect 31435 14028 32864 14056
rect 31435 14025 31447 14028
rect 31389 14019 31447 14025
rect 32858 14016 32864 14028
rect 32916 14016 32922 14068
rect 32953 14059 33011 14065
rect 32953 14025 32965 14059
rect 32999 14056 33011 14059
rect 34238 14056 34244 14068
rect 32999 14028 34244 14056
rect 32999 14025 33011 14028
rect 32953 14019 33011 14025
rect 34238 14016 34244 14028
rect 34296 14016 34302 14068
rect 35710 14016 35716 14068
rect 35768 14056 35774 14068
rect 35897 14059 35955 14065
rect 35897 14056 35909 14059
rect 35768 14028 35909 14056
rect 35768 14016 35774 14028
rect 35897 14025 35909 14028
rect 35943 14025 35955 14059
rect 35897 14019 35955 14025
rect 30834 13948 30840 14000
rect 30892 13988 30898 14000
rect 32493 13991 32551 13997
rect 32493 13988 32505 13991
rect 30892 13960 32505 13988
rect 30892 13948 30898 13960
rect 32493 13957 32505 13960
rect 32539 13957 32551 13991
rect 32493 13951 32551 13957
rect 32582 13948 32588 14000
rect 32640 13988 32646 14000
rect 32640 13960 33824 13988
rect 32640 13948 32646 13960
rect 29086 13920 29092 13932
rect 29047 13892 29092 13920
rect 29086 13880 29092 13892
rect 29144 13880 29150 13932
rect 29914 13920 29920 13932
rect 29875 13892 29920 13920
rect 29914 13880 29920 13892
rect 29972 13880 29978 13932
rect 30742 13880 30748 13932
rect 30800 13920 30806 13932
rect 31573 13923 31631 13929
rect 31573 13920 31585 13923
rect 30800 13892 31585 13920
rect 30800 13880 30806 13892
rect 31573 13889 31585 13892
rect 31619 13889 31631 13923
rect 31573 13883 31631 13889
rect 31662 13880 31668 13932
rect 31720 13920 31726 13932
rect 32125 13923 32183 13929
rect 32125 13920 32137 13923
rect 31720 13892 32137 13920
rect 31720 13880 31726 13892
rect 32125 13889 32137 13892
rect 32171 13889 32183 13923
rect 32125 13883 32183 13889
rect 32309 13923 32367 13929
rect 32309 13889 32321 13923
rect 32355 13920 32367 13923
rect 32674 13920 32680 13932
rect 32355 13892 32680 13920
rect 32355 13889 32367 13892
rect 32309 13883 32367 13889
rect 32674 13880 32680 13892
rect 32732 13880 32738 13932
rect 33134 13920 33140 13932
rect 33095 13892 33140 13920
rect 33134 13880 33140 13892
rect 33192 13880 33198 13932
rect 33796 13929 33824 13960
rect 33781 13923 33839 13929
rect 33781 13889 33793 13923
rect 33827 13889 33839 13923
rect 33781 13883 33839 13889
rect 34422 13880 34428 13932
rect 34480 13920 34486 13932
rect 34517 13923 34575 13929
rect 34517 13920 34529 13923
rect 34480 13892 34529 13920
rect 34480 13880 34486 13892
rect 34517 13889 34529 13892
rect 34563 13889 34575 13923
rect 34517 13883 34575 13889
rect 34606 13880 34612 13932
rect 34664 13920 34670 13932
rect 34773 13923 34831 13929
rect 34773 13920 34785 13923
rect 34664 13892 34785 13920
rect 34664 13880 34670 13892
rect 34773 13889 34785 13892
rect 34819 13889 34831 13923
rect 34773 13883 34831 13889
rect 34146 13852 34152 13864
rect 33612 13824 34152 13852
rect 33612 13793 33640 13824
rect 34146 13812 34152 13824
rect 34204 13812 34210 13864
rect 33597 13787 33655 13793
rect 33597 13753 33609 13787
rect 33643 13753 33655 13787
rect 33597 13747 33655 13753
rect 29181 13719 29239 13725
rect 29181 13716 29193 13719
rect 28966 13688 29193 13716
rect 29181 13685 29193 13688
rect 29227 13716 29239 13719
rect 34698 13716 34704 13728
rect 29227 13688 34704 13716
rect 29227 13685 29239 13688
rect 29181 13679 29239 13685
rect 34698 13676 34704 13688
rect 34756 13676 34762 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 5442 13472 5448 13524
rect 5500 13512 5506 13524
rect 6273 13515 6331 13521
rect 6273 13512 6285 13515
rect 5500 13484 6285 13512
rect 5500 13472 5506 13484
rect 6273 13481 6285 13484
rect 6319 13481 6331 13515
rect 6273 13475 6331 13481
rect 9122 13472 9128 13524
rect 9180 13512 9186 13524
rect 9309 13515 9367 13521
rect 9309 13512 9321 13515
rect 9180 13484 9321 13512
rect 9180 13472 9186 13484
rect 9309 13481 9321 13484
rect 9355 13481 9367 13515
rect 13630 13512 13636 13524
rect 9309 13475 9367 13481
rect 11440 13484 13636 13512
rect 8389 13447 8447 13453
rect 8389 13413 8401 13447
rect 8435 13444 8447 13447
rect 9214 13444 9220 13456
rect 8435 13416 9220 13444
rect 8435 13413 8447 13416
rect 8389 13407 8447 13413
rect 9214 13404 9220 13416
rect 9272 13404 9278 13456
rect 6454 13308 6460 13320
rect 6415 13280 6460 13308
rect 6454 13268 6460 13280
rect 6512 13268 6518 13320
rect 6822 13268 6828 13320
rect 6880 13308 6886 13320
rect 7009 13311 7067 13317
rect 7009 13308 7021 13311
rect 6880 13280 7021 13308
rect 6880 13268 6886 13280
rect 7009 13277 7021 13280
rect 7055 13308 7067 13311
rect 10045 13311 10103 13317
rect 10045 13308 10057 13311
rect 7055 13280 10057 13308
rect 7055 13277 7067 13280
rect 7009 13271 7067 13277
rect 10045 13277 10057 13280
rect 10091 13277 10103 13311
rect 10045 13271 10103 13277
rect 7276 13243 7334 13249
rect 7276 13209 7288 13243
rect 7322 13240 7334 13243
rect 7926 13240 7932 13252
rect 7322 13212 7932 13240
rect 7322 13209 7334 13212
rect 7276 13203 7334 13209
rect 7926 13200 7932 13212
rect 7984 13200 7990 13252
rect 8846 13200 8852 13252
rect 8904 13240 8910 13252
rect 8941 13243 8999 13249
rect 8941 13240 8953 13243
rect 8904 13212 8953 13240
rect 8904 13200 8910 13212
rect 8941 13209 8953 13212
rect 8987 13209 8999 13243
rect 9122 13240 9128 13252
rect 9083 13212 9128 13240
rect 8941 13203 8999 13209
rect 9122 13200 9128 13212
rect 9180 13200 9186 13252
rect 10318 13249 10324 13252
rect 10312 13203 10324 13249
rect 10376 13240 10382 13252
rect 10376 13212 10412 13240
rect 10318 13200 10324 13203
rect 10376 13200 10382 13212
rect 10226 13132 10232 13184
rect 10284 13172 10290 13184
rect 11440 13181 11468 13484
rect 13630 13472 13636 13484
rect 13688 13472 13694 13524
rect 14185 13515 14243 13521
rect 14185 13481 14197 13515
rect 14231 13512 14243 13515
rect 15194 13512 15200 13524
rect 14231 13484 15200 13512
rect 14231 13481 14243 13484
rect 14185 13475 14243 13481
rect 15194 13472 15200 13484
rect 15252 13472 15258 13524
rect 16942 13512 16948 13524
rect 15298 13484 16948 13512
rect 13449 13447 13507 13453
rect 13449 13413 13461 13447
rect 13495 13444 13507 13447
rect 14458 13444 14464 13456
rect 13495 13416 14464 13444
rect 13495 13413 13507 13416
rect 13449 13407 13507 13413
rect 14458 13404 14464 13416
rect 14516 13444 14522 13456
rect 15298 13444 15326 13484
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 17589 13515 17647 13521
rect 17589 13481 17601 13515
rect 17635 13512 17647 13515
rect 23658 13512 23664 13524
rect 17635 13484 19840 13512
rect 23619 13484 23664 13512
rect 17635 13481 17647 13484
rect 17589 13475 17647 13481
rect 14516 13416 15326 13444
rect 14516 13404 14522 13416
rect 16666 13404 16672 13456
rect 16724 13444 16730 13456
rect 17221 13447 17279 13453
rect 17221 13444 17233 13447
rect 16724 13416 17233 13444
rect 16724 13404 16730 13416
rect 17221 13413 17233 13416
rect 17267 13444 17279 13447
rect 17862 13444 17868 13456
rect 17267 13416 17868 13444
rect 17267 13413 17279 13416
rect 17221 13407 17279 13413
rect 17862 13404 17868 13416
rect 17920 13404 17926 13456
rect 18325 13447 18383 13453
rect 18325 13413 18337 13447
rect 18371 13413 18383 13447
rect 19334 13444 19340 13456
rect 18325 13407 18383 13413
rect 19260 13416 19340 13444
rect 12066 13376 12072 13388
rect 12027 13348 12072 13376
rect 12066 13336 12072 13348
rect 12124 13336 12130 13388
rect 13998 13336 14004 13388
rect 14056 13376 14062 13388
rect 17313 13379 17371 13385
rect 14056 13348 14320 13376
rect 14056 13336 14062 13348
rect 12084 13308 12112 13336
rect 12084 13280 14044 13308
rect 12336 13243 12394 13249
rect 12336 13209 12348 13243
rect 12382 13240 12394 13243
rect 12894 13240 12900 13252
rect 12382 13212 12900 13240
rect 12382 13209 12394 13212
rect 12336 13203 12394 13209
rect 12894 13200 12900 13212
rect 12952 13200 12958 13252
rect 14016 13240 14044 13280
rect 14090 13268 14096 13320
rect 14148 13308 14154 13320
rect 14292 13317 14320 13348
rect 17313 13345 17325 13379
rect 17359 13376 17371 13379
rect 17402 13376 17408 13388
rect 17359 13348 17408 13376
rect 17359 13345 17371 13348
rect 17313 13339 17371 13345
rect 17402 13336 17408 13348
rect 17460 13376 17466 13388
rect 18340 13376 18368 13407
rect 19260 13385 19288 13416
rect 19334 13404 19340 13416
rect 19392 13404 19398 13456
rect 19812 13444 19840 13484
rect 23658 13472 23664 13484
rect 23716 13472 23722 13524
rect 24486 13512 24492 13524
rect 24447 13484 24492 13512
rect 24486 13472 24492 13484
rect 24544 13512 24550 13524
rect 26418 13512 26424 13524
rect 24544 13484 26004 13512
rect 26331 13484 26424 13512
rect 24544 13472 24550 13484
rect 21542 13444 21548 13456
rect 19812 13416 21548 13444
rect 21542 13404 21548 13416
rect 21600 13404 21606 13456
rect 19245 13379 19303 13385
rect 19245 13376 19257 13379
rect 17460 13348 18368 13376
rect 19076 13348 19257 13376
rect 17460 13336 17466 13348
rect 14277 13311 14335 13317
rect 14148 13280 14193 13308
rect 14148 13268 14154 13280
rect 14277 13277 14289 13311
rect 14323 13277 14335 13311
rect 14277 13271 14335 13277
rect 15013 13311 15071 13317
rect 15013 13277 15025 13311
rect 15059 13308 15071 13311
rect 15102 13308 15108 13320
rect 15059 13280 15108 13308
rect 15059 13277 15071 13280
rect 15013 13271 15071 13277
rect 15102 13268 15108 13280
rect 15160 13268 15166 13320
rect 15470 13308 15476 13320
rect 15431 13280 15476 13308
rect 15470 13268 15476 13280
rect 15528 13268 15534 13320
rect 15562 13268 15568 13320
rect 15620 13308 15626 13320
rect 15930 13308 15936 13320
rect 15620 13280 15665 13308
rect 15891 13280 15936 13308
rect 15620 13268 15626 13280
rect 15930 13268 15936 13280
rect 15988 13268 15994 13320
rect 16758 13268 16764 13320
rect 16816 13308 16822 13320
rect 17126 13317 17132 13320
rect 16945 13311 17003 13317
rect 16945 13308 16957 13311
rect 16816 13280 16957 13308
rect 16816 13268 16822 13280
rect 16945 13277 16957 13280
rect 16991 13277 17003 13311
rect 16945 13271 17003 13277
rect 17092 13311 17132 13317
rect 17092 13277 17104 13311
rect 17092 13271 17132 13277
rect 17126 13268 17132 13271
rect 17184 13268 17190 13320
rect 17862 13268 17868 13320
rect 17920 13308 17926 13320
rect 18141 13311 18199 13317
rect 18141 13308 18153 13311
rect 17920 13280 18153 13308
rect 17920 13268 17926 13280
rect 18141 13277 18153 13280
rect 18187 13277 18199 13311
rect 18141 13271 18199 13277
rect 15286 13240 15292 13252
rect 14016 13212 15292 13240
rect 15286 13200 15292 13212
rect 15344 13240 15350 13252
rect 16114 13240 16120 13252
rect 15344 13212 16120 13240
rect 15344 13200 15350 13212
rect 16114 13200 16120 13212
rect 16172 13200 16178 13252
rect 16209 13243 16267 13249
rect 16209 13209 16221 13243
rect 16255 13240 16267 13243
rect 18782 13240 18788 13252
rect 16255 13212 18788 13240
rect 16255 13209 16267 13212
rect 16209 13203 16267 13209
rect 18782 13200 18788 13212
rect 18840 13200 18846 13252
rect 11425 13175 11483 13181
rect 11425 13172 11437 13175
rect 10284 13144 11437 13172
rect 10284 13132 10290 13144
rect 11425 13141 11437 13144
rect 11471 13141 11483 13175
rect 19076 13172 19104 13348
rect 19245 13345 19257 13348
rect 19291 13345 19303 13379
rect 19245 13339 19303 13345
rect 19705 13379 19763 13385
rect 19705 13345 19717 13379
rect 19751 13376 19763 13379
rect 20530 13376 20536 13388
rect 19751 13348 20536 13376
rect 19751 13345 19763 13348
rect 19705 13339 19763 13345
rect 20530 13336 20536 13348
rect 20588 13336 20594 13388
rect 24673 13379 24731 13385
rect 23676 13348 24624 13376
rect 19426 13308 19432 13320
rect 19387 13280 19432 13308
rect 19426 13268 19432 13280
rect 19484 13268 19490 13320
rect 23676 13317 23704 13348
rect 19797 13311 19855 13317
rect 19797 13277 19809 13311
rect 19843 13277 19855 13311
rect 19797 13271 19855 13277
rect 23661 13311 23719 13317
rect 23661 13277 23673 13311
rect 23707 13277 23719 13311
rect 23661 13271 23719 13277
rect 23845 13311 23903 13317
rect 23845 13277 23857 13311
rect 23891 13277 23903 13311
rect 24394 13308 24400 13320
rect 24355 13280 24400 13308
rect 23845 13271 23903 13277
rect 19150 13200 19156 13252
rect 19208 13240 19214 13252
rect 19812 13240 19840 13271
rect 19208 13212 19840 13240
rect 19208 13200 19214 13212
rect 23750 13200 23756 13252
rect 23808 13240 23814 13252
rect 23860 13240 23888 13271
rect 24394 13268 24400 13280
rect 24452 13268 24458 13320
rect 24596 13308 24624 13348
rect 24673 13345 24685 13379
rect 24719 13376 24731 13379
rect 24946 13376 24952 13388
rect 24719 13348 24952 13376
rect 24719 13345 24731 13348
rect 24673 13339 24731 13345
rect 24946 13336 24952 13348
rect 25004 13336 25010 13388
rect 25976 13376 26004 13484
rect 26418 13472 26424 13484
rect 26476 13512 26482 13524
rect 27154 13512 27160 13524
rect 26476 13484 27160 13512
rect 26476 13472 26482 13484
rect 27154 13472 27160 13484
rect 27212 13472 27218 13524
rect 27706 13512 27712 13524
rect 27667 13484 27712 13512
rect 27706 13472 27712 13484
rect 27764 13472 27770 13524
rect 30929 13515 30987 13521
rect 30929 13481 30941 13515
rect 30975 13512 30987 13515
rect 31662 13512 31668 13524
rect 30975 13484 31668 13512
rect 30975 13481 30987 13484
rect 30929 13475 30987 13481
rect 31662 13472 31668 13484
rect 31720 13472 31726 13524
rect 33413 13515 33471 13521
rect 33413 13481 33425 13515
rect 33459 13512 33471 13515
rect 34606 13512 34612 13524
rect 33459 13484 34612 13512
rect 33459 13481 33471 13484
rect 33413 13475 33471 13481
rect 34606 13472 34612 13484
rect 34664 13472 34670 13524
rect 35986 13512 35992 13524
rect 34716 13484 35992 13512
rect 26050 13404 26056 13456
rect 26108 13444 26114 13456
rect 32769 13447 32827 13453
rect 26108 13416 30604 13444
rect 26108 13404 26114 13416
rect 26329 13379 26387 13385
rect 26329 13376 26341 13379
rect 25976 13348 26341 13376
rect 26329 13345 26341 13348
rect 26375 13345 26387 13379
rect 26510 13376 26516 13388
rect 26471 13348 26516 13376
rect 26329 13339 26387 13345
rect 25038 13308 25044 13320
rect 24596 13280 25044 13308
rect 25038 13268 25044 13280
rect 25096 13308 25102 13320
rect 25593 13311 25651 13317
rect 25593 13308 25605 13311
rect 25096 13280 25605 13308
rect 25096 13268 25102 13280
rect 25593 13277 25605 13280
rect 25639 13277 25651 13311
rect 25593 13271 25651 13277
rect 25777 13311 25835 13317
rect 25777 13277 25789 13311
rect 25823 13277 25835 13311
rect 26234 13308 26240 13320
rect 26195 13280 26240 13308
rect 25777 13271 25835 13277
rect 24673 13243 24731 13249
rect 24673 13240 24685 13243
rect 23808 13212 24685 13240
rect 23808 13200 23814 13212
rect 24673 13209 24685 13212
rect 24719 13209 24731 13243
rect 25792 13240 25820 13271
rect 26234 13268 26240 13280
rect 26292 13268 26298 13320
rect 26344 13308 26372 13339
rect 26510 13336 26516 13348
rect 26568 13336 26574 13388
rect 27065 13379 27123 13385
rect 27065 13376 27077 13379
rect 26620 13348 27077 13376
rect 26620 13308 26648 13348
rect 27065 13345 27077 13348
rect 27111 13345 27123 13379
rect 27246 13376 27252 13388
rect 27207 13348 27252 13376
rect 27065 13339 27123 13345
rect 27246 13336 27252 13348
rect 27304 13336 27310 13388
rect 26970 13308 26976 13320
rect 26344 13280 26648 13308
rect 26931 13280 26976 13308
rect 26970 13268 26976 13280
rect 27028 13268 27034 13320
rect 27522 13268 27528 13320
rect 27580 13308 27586 13320
rect 27709 13311 27767 13317
rect 27709 13308 27721 13311
rect 27580 13280 27721 13308
rect 27580 13268 27586 13280
rect 27709 13277 27721 13280
rect 27755 13277 27767 13311
rect 27709 13271 27767 13277
rect 27893 13311 27951 13317
rect 27893 13277 27905 13311
rect 27939 13308 27951 13311
rect 28258 13308 28264 13320
rect 27939 13280 28264 13308
rect 27939 13277 27951 13280
rect 27893 13271 27951 13277
rect 28258 13268 28264 13280
rect 28316 13268 28322 13320
rect 30466 13308 30472 13320
rect 30427 13280 30472 13308
rect 30466 13268 30472 13280
rect 30524 13268 30530 13320
rect 30576 13308 30604 13416
rect 32769 13413 32781 13447
rect 32815 13444 32827 13447
rect 34716 13444 34744 13484
rect 35986 13472 35992 13484
rect 36044 13472 36050 13524
rect 32815 13416 34744 13444
rect 32815 13413 32827 13416
rect 32769 13407 32827 13413
rect 31113 13311 31171 13317
rect 31113 13308 31125 13311
rect 30576 13280 31125 13308
rect 31113 13277 31125 13280
rect 31159 13308 31171 13311
rect 31757 13311 31815 13317
rect 31757 13308 31769 13311
rect 31159 13280 31769 13308
rect 31159 13277 31171 13280
rect 31113 13271 31171 13277
rect 31757 13277 31769 13280
rect 31803 13308 31815 13311
rect 31846 13308 31852 13320
rect 31803 13280 31852 13308
rect 31803 13277 31815 13280
rect 31757 13271 31815 13277
rect 31846 13268 31852 13280
rect 31904 13268 31910 13320
rect 32953 13311 33011 13317
rect 32953 13277 32965 13311
rect 32999 13308 33011 13311
rect 33318 13308 33324 13320
rect 32999 13280 33324 13308
rect 32999 13277 33011 13280
rect 32953 13271 33011 13277
rect 33318 13268 33324 13280
rect 33376 13268 33382 13320
rect 33594 13308 33600 13320
rect 33555 13280 33600 13308
rect 33594 13268 33600 13280
rect 33652 13268 33658 13320
rect 34146 13268 34152 13320
rect 34204 13308 34210 13320
rect 34701 13311 34759 13317
rect 34701 13308 34713 13311
rect 34204 13280 34713 13308
rect 34204 13268 34210 13280
rect 34701 13277 34713 13280
rect 34747 13277 34759 13311
rect 34701 13271 34759 13277
rect 26878 13240 26884 13252
rect 25792 13212 26884 13240
rect 24673 13203 24731 13209
rect 26878 13200 26884 13212
rect 26936 13240 26942 13252
rect 27249 13243 27307 13249
rect 27249 13240 27261 13243
rect 26936 13212 27261 13240
rect 26936 13200 26942 13212
rect 27249 13209 27261 13212
rect 27295 13209 27307 13243
rect 27249 13203 27307 13209
rect 32858 13200 32864 13252
rect 32916 13240 32922 13252
rect 34946 13243 35004 13249
rect 34946 13240 34958 13243
rect 32916 13212 34958 13240
rect 32916 13200 32922 13212
rect 34946 13209 34958 13212
rect 34992 13209 35004 13243
rect 34946 13203 35004 13209
rect 19426 13172 19432 13184
rect 19076 13144 19432 13172
rect 11425 13135 11483 13141
rect 19426 13132 19432 13144
rect 19484 13132 19490 13184
rect 25682 13172 25688 13184
rect 25643 13144 25688 13172
rect 25682 13132 25688 13144
rect 25740 13132 25746 13184
rect 30282 13172 30288 13184
rect 30243 13144 30288 13172
rect 30282 13132 30288 13144
rect 30340 13132 30346 13184
rect 31573 13175 31631 13181
rect 31573 13141 31585 13175
rect 31619 13172 31631 13175
rect 32766 13172 32772 13184
rect 31619 13144 32772 13172
rect 31619 13141 31631 13144
rect 31573 13135 31631 13141
rect 32766 13132 32772 13144
rect 32824 13132 32830 13184
rect 33686 13132 33692 13184
rect 33744 13172 33750 13184
rect 36081 13175 36139 13181
rect 36081 13172 36093 13175
rect 33744 13144 36093 13172
rect 33744 13132 33750 13144
rect 36081 13141 36093 13144
rect 36127 13141 36139 13175
rect 36081 13135 36139 13141
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 4065 12971 4123 12977
rect 4065 12937 4077 12971
rect 4111 12968 4123 12971
rect 6086 12968 6092 12980
rect 4111 12940 6092 12968
rect 4111 12937 4123 12940
rect 4065 12931 4123 12937
rect 6086 12928 6092 12940
rect 6144 12928 6150 12980
rect 8386 12928 8392 12980
rect 8444 12968 8450 12980
rect 9030 12968 9036 12980
rect 8444 12940 9036 12968
rect 8444 12928 8450 12940
rect 9030 12928 9036 12940
rect 9088 12968 9094 12980
rect 9401 12971 9459 12977
rect 9401 12968 9413 12971
rect 9088 12940 9413 12968
rect 9088 12928 9094 12940
rect 9401 12937 9413 12940
rect 9447 12937 9459 12971
rect 20073 12971 20131 12977
rect 20073 12968 20085 12971
rect 9401 12931 9459 12937
rect 12406 12940 20085 12968
rect 2952 12903 3010 12909
rect 2952 12869 2964 12903
rect 2998 12900 3010 12903
rect 3694 12900 3700 12912
rect 2998 12872 3700 12900
rect 2998 12869 3010 12872
rect 2952 12863 3010 12869
rect 3694 12860 3700 12872
rect 3752 12860 3758 12912
rect 7644 12903 7702 12909
rect 7644 12869 7656 12903
rect 7690 12900 7702 12903
rect 8938 12900 8944 12912
rect 7690 12872 8944 12900
rect 7690 12869 7702 12872
rect 7644 12863 7702 12869
rect 8938 12860 8944 12872
rect 8996 12860 9002 12912
rect 9309 12903 9367 12909
rect 9309 12869 9321 12903
rect 9355 12900 9367 12903
rect 12406 12900 12434 12940
rect 20073 12937 20085 12940
rect 20119 12937 20131 12971
rect 20073 12931 20131 12937
rect 12894 12900 12900 12912
rect 9355 12872 12434 12900
rect 12855 12872 12900 12900
rect 9355 12869 9367 12872
rect 9309 12863 9367 12869
rect 12894 12860 12900 12872
rect 12952 12860 12958 12912
rect 14090 12860 14096 12912
rect 14148 12900 14154 12912
rect 14148 12872 15240 12900
rect 14148 12860 14154 12872
rect 15212 12844 15240 12872
rect 16390 12860 16396 12912
rect 16448 12900 16454 12912
rect 17034 12900 17040 12912
rect 16448 12872 17040 12900
rect 16448 12860 16454 12872
rect 17034 12860 17040 12872
rect 17092 12860 17098 12912
rect 17405 12903 17463 12909
rect 17405 12869 17417 12903
rect 17451 12900 17463 12903
rect 17586 12900 17592 12912
rect 17451 12872 17592 12900
rect 17451 12869 17463 12872
rect 17405 12863 17463 12869
rect 17586 12860 17592 12872
rect 17644 12860 17650 12912
rect 17678 12860 17684 12912
rect 17736 12900 17742 12912
rect 18141 12903 18199 12909
rect 18141 12900 18153 12903
rect 17736 12872 18153 12900
rect 17736 12860 17742 12872
rect 18141 12869 18153 12872
rect 18187 12869 18199 12903
rect 18141 12863 18199 12869
rect 19334 12860 19340 12912
rect 19392 12900 19398 12912
rect 19978 12900 19984 12912
rect 19392 12872 19437 12900
rect 19939 12872 19984 12900
rect 19392 12860 19398 12872
rect 19978 12860 19984 12872
rect 20036 12860 20042 12912
rect 20088 12900 20116 12931
rect 30184 12903 30242 12909
rect 20088 12872 21404 12900
rect 2682 12832 2688 12844
rect 2643 12804 2688 12832
rect 2682 12792 2688 12804
rect 2740 12792 2746 12844
rect 6822 12792 6828 12844
rect 6880 12832 6886 12844
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 6880 12804 7389 12832
rect 6880 12792 6886 12804
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 10413 12835 10471 12841
rect 10413 12832 10425 12835
rect 7377 12795 7435 12801
rect 7484 12804 10425 12832
rect 5258 12724 5264 12776
rect 5316 12764 5322 12776
rect 7484 12764 7512 12804
rect 10413 12801 10425 12804
rect 10459 12801 10471 12835
rect 10413 12795 10471 12801
rect 12802 12792 12808 12844
rect 12860 12832 12866 12844
rect 12989 12835 13047 12841
rect 12860 12804 12905 12832
rect 12860 12792 12866 12804
rect 12989 12801 13001 12835
rect 13035 12832 13047 12835
rect 13262 12832 13268 12844
rect 13035 12804 13268 12832
rect 13035 12801 13047 12804
rect 12989 12795 13047 12801
rect 10042 12764 10048 12776
rect 5316 12736 7512 12764
rect 10003 12736 10048 12764
rect 5316 12724 5322 12736
rect 10042 12724 10048 12736
rect 10100 12724 10106 12776
rect 10226 12764 10232 12776
rect 10187 12736 10232 12764
rect 10226 12724 10232 12736
rect 10284 12724 10290 12776
rect 10686 12724 10692 12776
rect 10744 12764 10750 12776
rect 11517 12767 11575 12773
rect 11517 12764 11529 12767
rect 10744 12736 11529 12764
rect 10744 12724 10750 12736
rect 11517 12733 11529 12736
rect 11563 12733 11575 12767
rect 11790 12764 11796 12776
rect 11751 12736 11796 12764
rect 11517 12727 11575 12733
rect 8757 12699 8815 12705
rect 8757 12665 8769 12699
rect 8803 12696 8815 12699
rect 9122 12696 9128 12708
rect 8803 12668 9128 12696
rect 8803 12665 8815 12668
rect 8757 12659 8815 12665
rect 9122 12656 9128 12668
rect 9180 12656 9186 12708
rect 10321 12699 10379 12705
rect 10321 12665 10333 12699
rect 10367 12696 10379 12699
rect 10410 12696 10416 12708
rect 10367 12668 10416 12696
rect 10367 12665 10379 12668
rect 10321 12659 10379 12665
rect 10410 12656 10416 12668
rect 10468 12696 10474 12708
rect 10870 12696 10876 12708
rect 10468 12668 10876 12696
rect 10468 12656 10474 12668
rect 10870 12656 10876 12668
rect 10928 12656 10934 12708
rect 10226 12628 10232 12640
rect 10187 12600 10232 12628
rect 10226 12588 10232 12600
rect 10284 12588 10290 12640
rect 11532 12628 11560 12727
rect 11790 12724 11796 12736
rect 11848 12724 11854 12776
rect 11808 12696 11836 12724
rect 13096 12696 13124 12804
rect 13262 12792 13268 12804
rect 13320 12792 13326 12844
rect 13998 12792 14004 12844
rect 14056 12832 14062 12844
rect 14921 12835 14979 12841
rect 14921 12832 14933 12835
rect 14056 12804 14933 12832
rect 14056 12792 14062 12804
rect 14921 12801 14933 12804
rect 14967 12801 14979 12835
rect 15194 12832 15200 12844
rect 15107 12804 15200 12832
rect 14921 12795 14979 12801
rect 15194 12792 15200 12804
rect 15252 12792 15258 12844
rect 16666 12832 16672 12844
rect 16627 12804 16672 12832
rect 16666 12792 16672 12804
rect 16724 12792 16730 12844
rect 16945 12835 17003 12841
rect 16945 12801 16957 12835
rect 16991 12801 17003 12835
rect 16945 12795 17003 12801
rect 11808 12668 13124 12696
rect 15212 12736 16344 12764
rect 15212 12628 15240 12736
rect 15473 12699 15531 12705
rect 15473 12665 15485 12699
rect 15519 12696 15531 12699
rect 15930 12696 15936 12708
rect 15519 12668 15936 12696
rect 15519 12665 15531 12668
rect 15473 12659 15531 12665
rect 15930 12656 15936 12668
rect 15988 12656 15994 12708
rect 16316 12696 16344 12736
rect 16390 12724 16396 12776
rect 16448 12764 16454 12776
rect 16960 12764 16988 12795
rect 16448 12736 16988 12764
rect 17604 12764 17632 12860
rect 18046 12832 18052 12844
rect 18007 12804 18052 12832
rect 18046 12792 18052 12804
rect 18104 12792 18110 12844
rect 18233 12835 18291 12841
rect 18233 12801 18245 12835
rect 18279 12801 18291 12835
rect 18233 12795 18291 12801
rect 18248 12764 18276 12795
rect 18322 12792 18328 12844
rect 18380 12832 18386 12844
rect 18417 12835 18475 12841
rect 18417 12832 18429 12835
rect 18380 12804 18429 12832
rect 18380 12792 18386 12804
rect 18417 12801 18429 12804
rect 18463 12801 18475 12835
rect 18417 12795 18475 12801
rect 18509 12835 18567 12841
rect 18509 12801 18521 12835
rect 18555 12832 18567 12835
rect 18598 12832 18604 12844
rect 18555 12804 18604 12832
rect 18555 12801 18567 12804
rect 18509 12795 18567 12801
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 18874 12792 18880 12844
rect 18932 12832 18938 12844
rect 19150 12832 19156 12844
rect 18932 12804 19156 12832
rect 18932 12792 18938 12804
rect 19150 12792 19156 12804
rect 19208 12792 19214 12844
rect 19426 12832 19432 12844
rect 19387 12804 19432 12832
rect 19426 12792 19432 12804
rect 19484 12792 19490 12844
rect 20530 12792 20536 12844
rect 20588 12832 20594 12844
rect 20625 12835 20683 12841
rect 20625 12832 20637 12835
rect 20588 12804 20637 12832
rect 20588 12792 20594 12804
rect 20625 12801 20637 12804
rect 20671 12801 20683 12835
rect 20625 12795 20683 12801
rect 20809 12835 20867 12841
rect 20809 12801 20821 12835
rect 20855 12832 20867 12835
rect 21266 12832 21272 12844
rect 20855 12804 21272 12832
rect 20855 12801 20867 12804
rect 20809 12795 20867 12801
rect 21266 12792 21272 12804
rect 21324 12792 21330 12844
rect 17604 12736 18276 12764
rect 18969 12767 19027 12773
rect 16448 12724 16454 12736
rect 18969 12733 18981 12767
rect 19015 12764 19027 12767
rect 19015 12736 21312 12764
rect 19015 12733 19027 12736
rect 18969 12727 19027 12733
rect 16758 12696 16764 12708
rect 16316 12668 16620 12696
rect 16719 12668 16764 12696
rect 11532 12600 15240 12628
rect 15289 12631 15347 12637
rect 15289 12597 15301 12631
rect 15335 12628 15347 12631
rect 15654 12628 15660 12640
rect 15335 12600 15660 12628
rect 15335 12597 15347 12600
rect 15289 12591 15347 12597
rect 15654 12588 15660 12600
rect 15712 12628 15718 12640
rect 16390 12628 16396 12640
rect 15712 12600 16396 12628
rect 15712 12588 15718 12600
rect 16390 12588 16396 12600
rect 16448 12588 16454 12640
rect 16592 12628 16620 12668
rect 16758 12656 16764 12668
rect 16816 12656 16822 12708
rect 17865 12699 17923 12705
rect 17865 12665 17877 12699
rect 17911 12696 17923 12699
rect 19426 12696 19432 12708
rect 17911 12668 19432 12696
rect 17911 12665 17923 12668
rect 17865 12659 17923 12665
rect 19426 12656 19432 12668
rect 19484 12656 19490 12708
rect 20898 12696 20904 12708
rect 20548 12668 20904 12696
rect 20548 12628 20576 12668
rect 20898 12656 20904 12668
rect 20956 12656 20962 12708
rect 20714 12628 20720 12640
rect 16592 12600 20576 12628
rect 20675 12600 20720 12628
rect 20714 12588 20720 12600
rect 20772 12588 20778 12640
rect 21284 12628 21312 12736
rect 21376 12696 21404 12872
rect 30184 12869 30196 12903
rect 30230 12900 30242 12903
rect 30282 12900 30288 12912
rect 30230 12872 30288 12900
rect 30230 12869 30242 12872
rect 30184 12863 30242 12869
rect 30282 12860 30288 12872
rect 30340 12860 30346 12912
rect 31662 12860 31668 12912
rect 31720 12900 31726 12912
rect 32585 12903 32643 12909
rect 32585 12900 32597 12903
rect 31720 12872 32597 12900
rect 31720 12860 31726 12872
rect 32585 12869 32597 12872
rect 32631 12869 32643 12903
rect 32585 12863 32643 12869
rect 23661 12835 23719 12841
rect 23661 12801 23673 12835
rect 23707 12832 23719 12835
rect 23750 12832 23756 12844
rect 23707 12804 23756 12832
rect 23707 12801 23719 12804
rect 23661 12795 23719 12801
rect 23750 12792 23756 12804
rect 23808 12792 23814 12844
rect 23845 12835 23903 12841
rect 23845 12801 23857 12835
rect 23891 12832 23903 12835
rect 25130 12832 25136 12844
rect 23891 12804 25136 12832
rect 23891 12801 23903 12804
rect 23845 12795 23903 12801
rect 25130 12792 25136 12804
rect 25188 12792 25194 12844
rect 28258 12832 28264 12844
rect 28219 12804 28264 12832
rect 28258 12792 28264 12804
rect 28316 12792 28322 12844
rect 28442 12832 28448 12844
rect 28403 12804 28448 12832
rect 28442 12792 28448 12804
rect 28500 12792 28506 12844
rect 28902 12832 28908 12844
rect 28863 12804 28908 12832
rect 28902 12792 28908 12804
rect 28960 12792 28966 12844
rect 29089 12835 29147 12841
rect 29089 12801 29101 12835
rect 29135 12801 29147 12835
rect 29089 12795 29147 12801
rect 32769 12835 32827 12841
rect 32769 12801 32781 12835
rect 32815 12832 32827 12835
rect 34054 12832 34060 12844
rect 32815 12804 34060 12832
rect 32815 12801 32827 12804
rect 32769 12795 32827 12801
rect 28350 12724 28356 12776
rect 28408 12764 28414 12776
rect 29104 12764 29132 12795
rect 34054 12792 34060 12804
rect 34112 12792 34118 12844
rect 29638 12764 29644 12776
rect 28408 12736 29644 12764
rect 28408 12724 28414 12736
rect 29638 12724 29644 12736
rect 29696 12724 29702 12776
rect 29914 12764 29920 12776
rect 29875 12736 29920 12764
rect 29914 12724 29920 12736
rect 29972 12724 29978 12776
rect 29086 12696 29092 12708
rect 21376 12668 29092 12696
rect 29086 12656 29092 12668
rect 29144 12656 29150 12708
rect 23474 12628 23480 12640
rect 21284 12600 23480 12628
rect 23474 12588 23480 12600
rect 23532 12588 23538 12640
rect 23658 12628 23664 12640
rect 23619 12600 23664 12628
rect 23658 12588 23664 12600
rect 23716 12588 23722 12640
rect 28166 12588 28172 12640
rect 28224 12628 28230 12640
rect 28261 12631 28319 12637
rect 28261 12628 28273 12631
rect 28224 12600 28273 12628
rect 28224 12588 28230 12600
rect 28261 12597 28273 12600
rect 28307 12597 28319 12631
rect 28261 12591 28319 12597
rect 28718 12588 28724 12640
rect 28776 12628 28782 12640
rect 28905 12631 28963 12637
rect 28905 12628 28917 12631
rect 28776 12600 28917 12628
rect 28776 12588 28782 12600
rect 28905 12597 28917 12600
rect 28951 12597 28963 12631
rect 31294 12628 31300 12640
rect 31255 12600 31300 12628
rect 28905 12591 28963 12597
rect 31294 12588 31300 12600
rect 31352 12588 31358 12640
rect 31754 12588 31760 12640
rect 31812 12628 31818 12640
rect 32953 12631 33011 12637
rect 32953 12628 32965 12631
rect 31812 12600 32965 12628
rect 31812 12588 31818 12600
rect 32953 12597 32965 12600
rect 32999 12597 33011 12631
rect 32953 12591 33011 12597
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 8294 12384 8300 12436
rect 8352 12424 8358 12436
rect 8389 12427 8447 12433
rect 8389 12424 8401 12427
rect 8352 12396 8401 12424
rect 8352 12384 8358 12396
rect 8389 12393 8401 12396
rect 8435 12393 8447 12427
rect 10318 12424 10324 12436
rect 10279 12396 10324 12424
rect 8389 12387 8447 12393
rect 10318 12384 10324 12396
rect 10376 12384 10382 12436
rect 14274 12424 14280 12436
rect 14235 12396 14280 12424
rect 14274 12384 14280 12396
rect 14332 12384 14338 12436
rect 14369 12427 14427 12433
rect 14369 12393 14381 12427
rect 14415 12424 14427 12427
rect 15746 12424 15752 12436
rect 14415 12396 15752 12424
rect 14415 12393 14427 12396
rect 14369 12387 14427 12393
rect 15746 12384 15752 12396
rect 15804 12384 15810 12436
rect 16301 12427 16359 12433
rect 16301 12393 16313 12427
rect 16347 12424 16359 12427
rect 16390 12424 16396 12436
rect 16347 12396 16396 12424
rect 16347 12393 16359 12396
rect 16301 12387 16359 12393
rect 16390 12384 16396 12396
rect 16448 12384 16454 12436
rect 16758 12384 16764 12436
rect 16816 12424 16822 12436
rect 17497 12427 17555 12433
rect 16816 12396 17448 12424
rect 16816 12384 16822 12396
rect 14458 12356 14464 12368
rect 14292 12328 14464 12356
rect 6822 12248 6828 12300
rect 6880 12288 6886 12300
rect 14292 12297 14320 12328
rect 14458 12316 14464 12328
rect 14516 12316 14522 12368
rect 15657 12359 15715 12365
rect 15657 12325 15669 12359
rect 15703 12356 15715 12359
rect 16850 12356 16856 12368
rect 15703 12328 16856 12356
rect 15703 12325 15715 12328
rect 15657 12319 15715 12325
rect 16850 12316 16856 12328
rect 16908 12356 16914 12368
rect 16991 12359 17049 12365
rect 16991 12356 17003 12359
rect 16908 12328 17003 12356
rect 16908 12316 16914 12328
rect 16991 12325 17003 12328
rect 17037 12325 17049 12359
rect 16991 12319 17049 12325
rect 17129 12359 17187 12365
rect 17129 12325 17141 12359
rect 17175 12325 17187 12359
rect 17420 12356 17448 12396
rect 17497 12393 17509 12427
rect 17543 12424 17555 12427
rect 17678 12424 17684 12436
rect 17543 12396 17684 12424
rect 17543 12393 17555 12396
rect 17497 12387 17555 12393
rect 17678 12384 17684 12396
rect 17736 12384 17742 12436
rect 19794 12424 19800 12436
rect 19755 12396 19800 12424
rect 19794 12384 19800 12396
rect 19852 12384 19858 12436
rect 22925 12427 22983 12433
rect 22925 12393 22937 12427
rect 22971 12393 22983 12427
rect 22925 12387 22983 12393
rect 17862 12356 17868 12368
rect 17420 12328 17868 12356
rect 17129 12319 17187 12325
rect 7009 12291 7067 12297
rect 7009 12288 7021 12291
rect 6880 12260 7021 12288
rect 6880 12248 6886 12260
rect 7009 12257 7021 12260
rect 7055 12257 7067 12291
rect 7009 12251 7067 12257
rect 14277 12291 14335 12297
rect 14277 12257 14289 12291
rect 14323 12257 14335 12291
rect 14277 12251 14335 12257
rect 15470 12248 15476 12300
rect 15528 12288 15534 12300
rect 16482 12288 16488 12300
rect 15528 12260 16488 12288
rect 15528 12248 15534 12260
rect 16482 12248 16488 12260
rect 16540 12288 16546 12300
rect 17144 12288 17172 12319
rect 17862 12316 17868 12328
rect 17920 12356 17926 12368
rect 18233 12359 18291 12365
rect 18233 12356 18245 12359
rect 17920 12328 18245 12356
rect 17920 12316 17926 12328
rect 18233 12325 18245 12328
rect 18279 12325 18291 12359
rect 22940 12356 22968 12387
rect 23474 12384 23480 12436
rect 23532 12424 23538 12436
rect 26970 12424 26976 12436
rect 23532 12396 26648 12424
rect 26931 12396 26976 12424
rect 23532 12384 23538 12396
rect 22940 12328 23612 12356
rect 18233 12319 18291 12325
rect 16540 12260 17172 12288
rect 17221 12291 17279 12297
rect 16540 12248 16546 12260
rect 17221 12257 17233 12291
rect 17267 12257 17279 12291
rect 17221 12251 17279 12257
rect 22925 12291 22983 12297
rect 22925 12257 22937 12291
rect 22971 12257 22983 12291
rect 22925 12251 22983 12257
rect 9766 12220 9772 12232
rect 9727 12192 9772 12220
rect 9766 12180 9772 12192
rect 9824 12180 9830 12232
rect 10226 12220 10232 12232
rect 10187 12192 10232 12220
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 10410 12220 10416 12232
rect 10371 12192 10416 12220
rect 10410 12180 10416 12192
rect 10468 12220 10474 12232
rect 11790 12220 11796 12232
rect 10468 12192 11796 12220
rect 10468 12180 10474 12192
rect 11790 12180 11796 12192
rect 11848 12180 11854 12232
rect 14461 12223 14519 12229
rect 14461 12189 14473 12223
rect 14507 12220 14519 12223
rect 15102 12220 15108 12232
rect 14507 12192 15108 12220
rect 14507 12189 14519 12192
rect 14461 12183 14519 12189
rect 15102 12180 15108 12192
rect 15160 12180 15166 12232
rect 15289 12223 15347 12229
rect 15289 12189 15301 12223
rect 15335 12220 15347 12223
rect 16022 12220 16028 12232
rect 15335 12192 16028 12220
rect 15335 12189 15347 12192
rect 15289 12183 15347 12189
rect 16022 12180 16028 12192
rect 16080 12220 16086 12232
rect 16117 12223 16175 12229
rect 16117 12220 16129 12223
rect 16080 12192 16129 12220
rect 16080 12180 16086 12192
rect 16117 12189 16129 12192
rect 16163 12189 16175 12223
rect 17236 12220 17264 12251
rect 17954 12220 17960 12232
rect 17236 12192 17960 12220
rect 16117 12183 16175 12189
rect 17954 12180 17960 12192
rect 18012 12220 18018 12232
rect 18049 12223 18107 12229
rect 18049 12220 18061 12223
rect 18012 12192 18061 12220
rect 18012 12180 18018 12192
rect 18049 12189 18061 12192
rect 18095 12189 18107 12223
rect 18049 12183 18107 12189
rect 19242 12180 19248 12232
rect 19300 12220 19306 12232
rect 20441 12223 20499 12229
rect 20441 12220 20453 12223
rect 19300 12192 20453 12220
rect 19300 12180 19306 12192
rect 20441 12189 20453 12192
rect 20487 12220 20499 12223
rect 21818 12220 21824 12232
rect 20487 12192 21824 12220
rect 20487 12189 20499 12192
rect 20441 12183 20499 12189
rect 21818 12180 21824 12192
rect 21876 12180 21882 12232
rect 7276 12155 7334 12161
rect 7276 12121 7288 12155
rect 7322 12152 7334 12155
rect 7322 12124 9628 12152
rect 7322 12121 7334 12124
rect 7276 12115 7334 12121
rect 9600 12093 9628 12124
rect 12158 12112 12164 12164
rect 12216 12152 12222 12164
rect 14090 12152 14096 12164
rect 12216 12124 14096 12152
rect 12216 12112 12222 12124
rect 14090 12112 14096 12124
rect 14148 12112 14154 12164
rect 15378 12112 15384 12164
rect 15436 12152 15442 12164
rect 15473 12155 15531 12161
rect 15473 12152 15485 12155
rect 15436 12124 15485 12152
rect 15436 12112 15442 12124
rect 15473 12121 15485 12124
rect 15519 12121 15531 12155
rect 15473 12115 15531 12121
rect 16390 12112 16396 12164
rect 16448 12152 16454 12164
rect 16853 12155 16911 12161
rect 16853 12152 16865 12155
rect 16448 12124 16865 12152
rect 16448 12112 16454 12124
rect 16853 12121 16865 12124
rect 16899 12121 16911 12155
rect 16853 12115 16911 12121
rect 18322 12112 18328 12164
rect 18380 12152 18386 12164
rect 20714 12161 20720 12164
rect 19705 12155 19763 12161
rect 19705 12152 19717 12155
rect 18380 12124 19717 12152
rect 18380 12112 18386 12124
rect 19705 12121 19717 12124
rect 19751 12121 19763 12155
rect 19705 12115 19763 12121
rect 20708 12115 20720 12161
rect 20772 12152 20778 12164
rect 22738 12152 22744 12164
rect 20772 12124 20808 12152
rect 22699 12124 22744 12152
rect 20714 12112 20720 12115
rect 20772 12112 20778 12124
rect 22738 12112 22744 12124
rect 22796 12112 22802 12164
rect 22940 12152 22968 12251
rect 23014 12248 23020 12300
rect 23072 12288 23078 12300
rect 23072 12260 23117 12288
rect 23072 12248 23078 12260
rect 23109 12223 23167 12229
rect 23109 12189 23121 12223
rect 23155 12220 23167 12223
rect 23474 12220 23480 12232
rect 23155 12192 23480 12220
rect 23155 12189 23167 12192
rect 23109 12183 23167 12189
rect 23474 12180 23480 12192
rect 23532 12180 23538 12232
rect 23584 12229 23612 12328
rect 26620 12288 26648 12396
rect 26970 12384 26976 12396
rect 27028 12384 27034 12436
rect 30466 12384 30472 12436
rect 30524 12424 30530 12436
rect 30929 12427 30987 12433
rect 30929 12424 30941 12427
rect 30524 12396 30941 12424
rect 30524 12384 30530 12396
rect 30929 12393 30941 12396
rect 30975 12393 30987 12427
rect 30929 12387 30987 12393
rect 32582 12384 32588 12436
rect 32640 12424 32646 12436
rect 34146 12424 34152 12436
rect 32640 12396 34152 12424
rect 32640 12384 32646 12396
rect 34146 12384 34152 12396
rect 34204 12384 34210 12436
rect 29549 12359 29607 12365
rect 29549 12325 29561 12359
rect 29595 12356 29607 12359
rect 35526 12356 35532 12368
rect 29595 12328 35532 12356
rect 29595 12325 29607 12328
rect 29549 12319 29607 12325
rect 35526 12316 35532 12328
rect 35584 12316 35590 12368
rect 27525 12291 27583 12297
rect 27525 12288 27537 12291
rect 26620 12260 27537 12288
rect 27525 12257 27537 12260
rect 27571 12288 27583 12291
rect 28350 12288 28356 12300
rect 27571 12260 28356 12288
rect 27571 12257 27583 12260
rect 27525 12251 27583 12257
rect 28350 12248 28356 12260
rect 28408 12248 28414 12300
rect 28460 12260 29040 12288
rect 28460 12232 28488 12260
rect 23569 12223 23627 12229
rect 23569 12189 23581 12223
rect 23615 12189 23627 12223
rect 23569 12183 23627 12189
rect 23753 12223 23811 12229
rect 23753 12189 23765 12223
rect 23799 12220 23811 12223
rect 24118 12220 24124 12232
rect 23799 12192 24124 12220
rect 23799 12189 23811 12192
rect 23753 12183 23811 12189
rect 24118 12180 24124 12192
rect 24176 12180 24182 12232
rect 24949 12223 25007 12229
rect 24949 12189 24961 12223
rect 24995 12189 25007 12223
rect 25130 12220 25136 12232
rect 25091 12192 25136 12220
rect 24949 12183 25007 12189
rect 24854 12152 24860 12164
rect 22940 12124 24860 12152
rect 24854 12112 24860 12124
rect 24912 12112 24918 12164
rect 24964 12152 24992 12183
rect 25130 12180 25136 12192
rect 25188 12180 25194 12232
rect 25590 12220 25596 12232
rect 25551 12192 25596 12220
rect 25590 12180 25596 12192
rect 25648 12180 25654 12232
rect 25682 12180 25688 12232
rect 25740 12220 25746 12232
rect 25849 12223 25907 12229
rect 25849 12220 25861 12223
rect 25740 12192 25861 12220
rect 25740 12180 25746 12192
rect 25849 12189 25861 12192
rect 25895 12189 25907 12223
rect 27798 12220 27804 12232
rect 27759 12192 27804 12220
rect 25849 12183 25907 12189
rect 27798 12180 27804 12192
rect 27856 12220 27862 12232
rect 28442 12220 28448 12232
rect 27856 12192 28448 12220
rect 27856 12180 27862 12192
rect 28442 12180 28448 12192
rect 28500 12180 28506 12232
rect 28810 12220 28816 12232
rect 28771 12192 28816 12220
rect 28810 12180 28816 12192
rect 28868 12180 28874 12232
rect 29012 12229 29040 12260
rect 32766 12248 32772 12300
rect 32824 12248 32830 12300
rect 28997 12223 29055 12229
rect 28997 12189 29009 12223
rect 29043 12189 29055 12223
rect 29546 12220 29552 12232
rect 29507 12192 29552 12220
rect 28997 12183 29055 12189
rect 29546 12180 29552 12192
rect 29604 12180 29610 12232
rect 29638 12180 29644 12232
rect 29696 12220 29702 12232
rect 29733 12223 29791 12229
rect 29733 12220 29745 12223
rect 29696 12192 29745 12220
rect 29696 12180 29702 12192
rect 29733 12189 29745 12192
rect 29779 12189 29791 12223
rect 29733 12183 29791 12189
rect 30745 12223 30803 12229
rect 30745 12189 30757 12223
rect 30791 12220 30803 12223
rect 31294 12220 31300 12232
rect 30791 12192 31300 12220
rect 30791 12189 30803 12192
rect 30745 12183 30803 12189
rect 31294 12180 31300 12192
rect 31352 12180 31358 12232
rect 31757 12223 31815 12229
rect 31757 12220 31769 12223
rect 31404 12192 31769 12220
rect 26418 12152 26424 12164
rect 24964 12124 26424 12152
rect 26418 12112 26424 12124
rect 26476 12112 26482 12164
rect 30561 12155 30619 12161
rect 30561 12121 30573 12155
rect 30607 12152 30619 12155
rect 31404 12152 31432 12192
rect 31757 12189 31769 12192
rect 31803 12220 31815 12223
rect 31846 12220 31852 12232
rect 31803 12192 31852 12220
rect 31803 12189 31815 12192
rect 31757 12183 31815 12189
rect 31846 12180 31852 12192
rect 31904 12180 31910 12232
rect 32784 12220 32812 12248
rect 33413 12223 33471 12229
rect 33413 12220 33425 12223
rect 32784 12192 33425 12220
rect 33413 12189 33425 12192
rect 33459 12189 33471 12223
rect 33413 12183 33471 12189
rect 32122 12152 32128 12164
rect 30607 12124 31432 12152
rect 31726 12124 32128 12152
rect 30607 12121 30619 12124
rect 30561 12115 30619 12121
rect 9585 12087 9643 12093
rect 9585 12053 9597 12087
rect 9631 12053 9643 12087
rect 9585 12047 9643 12053
rect 18966 12044 18972 12096
rect 19024 12084 19030 12096
rect 20070 12084 20076 12096
rect 19024 12056 20076 12084
rect 19024 12044 19030 12056
rect 20070 12044 20076 12056
rect 20128 12084 20134 12096
rect 21821 12087 21879 12093
rect 21821 12084 21833 12087
rect 20128 12056 21833 12084
rect 20128 12044 20134 12056
rect 21821 12053 21833 12056
rect 21867 12053 21879 12087
rect 21821 12047 21879 12053
rect 23753 12087 23811 12093
rect 23753 12053 23765 12087
rect 23799 12084 23811 12087
rect 24026 12084 24032 12096
rect 23799 12056 24032 12084
rect 23799 12053 23811 12056
rect 23753 12047 23811 12053
rect 24026 12044 24032 12056
rect 24084 12044 24090 12096
rect 25041 12087 25099 12093
rect 25041 12053 25053 12087
rect 25087 12084 25099 12087
rect 25958 12084 25964 12096
rect 25087 12056 25964 12084
rect 25087 12053 25099 12056
rect 25041 12047 25099 12053
rect 25958 12044 25964 12056
rect 26016 12044 26022 12096
rect 28905 12087 28963 12093
rect 28905 12053 28917 12087
rect 28951 12084 28963 12087
rect 30742 12084 30748 12096
rect 28951 12056 30748 12084
rect 28951 12053 28963 12056
rect 28905 12047 28963 12053
rect 30742 12044 30748 12056
rect 30800 12044 30806 12096
rect 31573 12087 31631 12093
rect 31573 12053 31585 12087
rect 31619 12084 31631 12087
rect 31726 12084 31754 12124
rect 32122 12112 32128 12124
rect 32180 12152 32186 12164
rect 32585 12155 32643 12161
rect 32585 12152 32597 12155
rect 32180 12124 32597 12152
rect 32180 12112 32186 12124
rect 32585 12121 32597 12124
rect 32631 12121 32643 12155
rect 32585 12115 32643 12121
rect 32769 12155 32827 12161
rect 32769 12121 32781 12155
rect 32815 12152 32827 12155
rect 33226 12152 33232 12164
rect 32815 12124 33232 12152
rect 32815 12121 32827 12124
rect 32769 12115 32827 12121
rect 33226 12112 33232 12124
rect 33284 12112 33290 12164
rect 33594 12152 33600 12164
rect 33555 12124 33600 12152
rect 33594 12112 33600 12124
rect 33652 12112 33658 12164
rect 31619 12056 31754 12084
rect 32953 12087 33011 12093
rect 31619 12053 31631 12056
rect 31573 12047 31631 12053
rect 32953 12053 32965 12087
rect 32999 12084 33011 12087
rect 33686 12084 33692 12096
rect 32999 12056 33692 12084
rect 32999 12053 33011 12056
rect 32953 12047 33011 12053
rect 33686 12044 33692 12056
rect 33744 12044 33750 12096
rect 33778 12044 33784 12096
rect 33836 12084 33842 12096
rect 33836 12056 33881 12084
rect 33836 12044 33842 12056
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 7926 11880 7932 11892
rect 7887 11852 7932 11880
rect 7926 11840 7932 11852
rect 7984 11840 7990 11892
rect 10870 11840 10876 11892
rect 10928 11880 10934 11892
rect 13541 11883 13599 11889
rect 13541 11880 13553 11883
rect 10928 11852 13553 11880
rect 10928 11840 10934 11852
rect 13541 11849 13553 11852
rect 13587 11849 13599 11883
rect 17126 11880 17132 11892
rect 13541 11843 13599 11849
rect 16868 11852 17132 11880
rect 16868 11824 16896 11852
rect 17126 11840 17132 11852
rect 17184 11840 17190 11892
rect 17313 11883 17371 11889
rect 17313 11849 17325 11883
rect 17359 11880 17371 11883
rect 18046 11880 18052 11892
rect 17359 11852 18052 11880
rect 17359 11849 17371 11852
rect 17313 11843 17371 11849
rect 18046 11840 18052 11852
rect 18104 11840 18110 11892
rect 19061 11883 19119 11889
rect 19061 11849 19073 11883
rect 19107 11880 19119 11883
rect 19978 11880 19984 11892
rect 19107 11852 19984 11880
rect 19107 11849 19119 11852
rect 19061 11843 19119 11849
rect 19978 11840 19984 11852
rect 20036 11840 20042 11892
rect 21358 11840 21364 11892
rect 21416 11880 21422 11892
rect 23201 11883 23259 11889
rect 23201 11880 23213 11883
rect 21416 11852 23213 11880
rect 21416 11840 21422 11852
rect 23201 11849 23213 11852
rect 23247 11849 23259 11883
rect 23201 11843 23259 11849
rect 24854 11840 24860 11892
rect 24912 11880 24918 11892
rect 25133 11883 25191 11889
rect 25133 11880 25145 11883
rect 24912 11852 25145 11880
rect 24912 11840 24918 11852
rect 25133 11849 25145 11852
rect 25179 11880 25191 11883
rect 25222 11880 25228 11892
rect 25179 11852 25228 11880
rect 25179 11849 25191 11852
rect 25133 11843 25191 11849
rect 25222 11840 25228 11852
rect 25280 11840 25286 11892
rect 28442 11840 28448 11892
rect 28500 11880 28506 11892
rect 28718 11880 28724 11892
rect 28500 11852 28724 11880
rect 28500 11840 28506 11852
rect 28718 11840 28724 11852
rect 28776 11840 28782 11892
rect 34054 11880 34060 11892
rect 34015 11852 34060 11880
rect 34054 11840 34060 11852
rect 34112 11840 34118 11892
rect 9214 11772 9220 11824
rect 9272 11812 9278 11824
rect 14369 11815 14427 11821
rect 14369 11812 14381 11815
rect 9272 11784 14381 11812
rect 9272 11772 9278 11784
rect 14369 11781 14381 11784
rect 14415 11781 14427 11815
rect 16850 11812 16856 11824
rect 16763 11784 16856 11812
rect 14369 11775 14427 11781
rect 16850 11772 16856 11784
rect 16908 11772 16914 11824
rect 19683 11815 19741 11821
rect 19683 11781 19695 11815
rect 19729 11812 19741 11815
rect 20530 11812 20536 11824
rect 19729 11784 20536 11812
rect 19729 11781 19741 11784
rect 19683 11775 19741 11781
rect 20530 11772 20536 11784
rect 20588 11772 20594 11824
rect 24026 11821 24032 11824
rect 24020 11812 24032 11821
rect 21836 11784 23796 11812
rect 23987 11784 24032 11812
rect 21836 11756 21864 11784
rect 8110 11744 8116 11756
rect 8071 11716 8116 11744
rect 8110 11704 8116 11716
rect 8168 11704 8174 11756
rect 12618 11744 12624 11756
rect 12579 11716 12624 11744
rect 12618 11704 12624 11716
rect 12676 11704 12682 11756
rect 13449 11747 13507 11753
rect 13449 11713 13461 11747
rect 13495 11744 13507 11747
rect 13538 11744 13544 11756
rect 13495 11716 13544 11744
rect 13495 11713 13507 11716
rect 13449 11707 13507 11713
rect 13538 11704 13544 11716
rect 13596 11704 13602 11756
rect 16758 11704 16764 11756
rect 16816 11744 16822 11756
rect 17129 11747 17187 11753
rect 17129 11744 17141 11747
rect 16816 11716 17141 11744
rect 16816 11704 16822 11716
rect 17129 11713 17141 11716
rect 17175 11713 17187 11747
rect 17129 11707 17187 11713
rect 18322 11704 18328 11756
rect 18380 11744 18386 11756
rect 18877 11747 18935 11753
rect 18877 11744 18889 11747
rect 18380 11716 18889 11744
rect 18380 11704 18386 11716
rect 18877 11713 18889 11716
rect 18923 11713 18935 11747
rect 18877 11707 18935 11713
rect 18966 11704 18972 11756
rect 19024 11744 19030 11756
rect 19981 11747 20039 11753
rect 19981 11744 19993 11747
rect 19024 11716 19993 11744
rect 19024 11704 19030 11716
rect 19981 11713 19993 11716
rect 20027 11713 20039 11747
rect 21082 11744 21088 11756
rect 21043 11716 21088 11744
rect 19981 11707 20039 11713
rect 21082 11704 21088 11716
rect 21140 11704 21146 11756
rect 21266 11744 21272 11756
rect 21227 11716 21272 11744
rect 21266 11704 21272 11716
rect 21324 11704 21330 11756
rect 21818 11744 21824 11756
rect 21779 11716 21824 11744
rect 21818 11704 21824 11716
rect 21876 11704 21882 11756
rect 23768 11753 23796 11784
rect 24020 11775 24032 11784
rect 24026 11772 24032 11775
rect 24084 11772 24090 11824
rect 24118 11772 24124 11824
rect 24176 11812 24182 11824
rect 24176 11784 25820 11812
rect 24176 11772 24182 11784
rect 22077 11747 22135 11753
rect 22077 11744 22089 11747
rect 21928 11716 22089 11744
rect 12894 11676 12900 11688
rect 12855 11648 12900 11676
rect 12894 11636 12900 11648
rect 12952 11636 12958 11688
rect 16114 11676 16120 11688
rect 16075 11648 16120 11676
rect 16114 11636 16120 11648
rect 16172 11636 16178 11688
rect 16390 11636 16396 11688
rect 16448 11676 16454 11688
rect 16945 11679 17003 11685
rect 16945 11676 16957 11679
rect 16448 11648 16957 11676
rect 16448 11636 16454 11648
rect 16945 11645 16957 11648
rect 16991 11645 17003 11679
rect 16945 11639 17003 11645
rect 19797 11679 19855 11685
rect 19797 11645 19809 11679
rect 19843 11676 19855 11679
rect 20070 11676 20076 11688
rect 19843 11648 20076 11676
rect 19843 11645 19855 11648
rect 19797 11639 19855 11645
rect 20070 11636 20076 11648
rect 20128 11636 20134 11688
rect 21177 11679 21235 11685
rect 21177 11645 21189 11679
rect 21223 11676 21235 11679
rect 21928 11676 21956 11716
rect 22077 11713 22089 11716
rect 22123 11713 22135 11747
rect 22077 11707 22135 11713
rect 23753 11747 23811 11753
rect 23753 11713 23765 11747
rect 23799 11713 23811 11747
rect 23753 11707 23811 11713
rect 24946 11704 24952 11756
rect 25004 11744 25010 11756
rect 25792 11753 25820 11784
rect 27614 11772 27620 11824
rect 27672 11812 27678 11824
rect 27672 11784 28580 11812
rect 27672 11772 27678 11784
rect 25593 11747 25651 11753
rect 25593 11744 25605 11747
rect 25004 11716 25605 11744
rect 25004 11704 25010 11716
rect 25593 11713 25605 11716
rect 25639 11713 25651 11747
rect 25593 11707 25651 11713
rect 25777 11747 25835 11753
rect 25777 11713 25789 11747
rect 25823 11713 25835 11747
rect 25777 11707 25835 11713
rect 26878 11704 26884 11756
rect 26936 11744 26942 11756
rect 26973 11747 27031 11753
rect 26973 11744 26985 11747
rect 26936 11716 26985 11744
rect 26936 11704 26942 11716
rect 26973 11713 26985 11716
rect 27019 11713 27031 11747
rect 26973 11707 27031 11713
rect 27157 11747 27215 11753
rect 27157 11713 27169 11747
rect 27203 11713 27215 11747
rect 28350 11744 28356 11756
rect 28311 11716 28356 11744
rect 27157 11707 27215 11713
rect 21223 11648 21956 11676
rect 21223 11645 21235 11648
rect 21177 11639 21235 11645
rect 25130 11636 25136 11688
rect 25188 11676 25194 11688
rect 27172 11676 27200 11707
rect 28350 11704 28356 11716
rect 28408 11704 28414 11756
rect 28552 11753 28580 11784
rect 28537 11747 28595 11753
rect 28537 11713 28549 11747
rect 28583 11713 28595 11747
rect 28537 11707 28595 11713
rect 31573 11747 31631 11753
rect 31573 11713 31585 11747
rect 31619 11744 31631 11747
rect 31754 11744 31760 11756
rect 31619 11716 31760 11744
rect 31619 11713 31631 11716
rect 31573 11707 31631 11713
rect 31754 11704 31760 11716
rect 31812 11704 31818 11756
rect 32933 11747 32991 11753
rect 32933 11744 32945 11747
rect 32324 11716 32945 11744
rect 27798 11676 27804 11688
rect 25188 11648 27804 11676
rect 25188 11636 25194 11648
rect 27798 11636 27804 11648
rect 27856 11636 27862 11688
rect 28718 11676 28724 11688
rect 28679 11648 28724 11676
rect 28718 11636 28724 11648
rect 28776 11636 28782 11688
rect 32324 11676 32352 11716
rect 32933 11713 32945 11716
rect 32979 11713 32991 11747
rect 32933 11707 32991 11713
rect 33686 11704 33692 11756
rect 33744 11744 33750 11756
rect 34701 11747 34759 11753
rect 34701 11744 34713 11747
rect 33744 11716 34713 11744
rect 33744 11704 33750 11716
rect 34701 11713 34713 11716
rect 34747 11713 34759 11747
rect 34701 11707 34759 11713
rect 31726 11648 32352 11676
rect 15746 11568 15752 11620
rect 15804 11608 15810 11620
rect 15804 11580 19334 11608
rect 15804 11568 15810 11580
rect 12342 11500 12348 11552
rect 12400 11540 12406 11552
rect 12437 11543 12495 11549
rect 12437 11540 12449 11543
rect 12400 11512 12449 11540
rect 12400 11500 12406 11512
rect 12437 11509 12449 11512
rect 12483 11509 12495 11543
rect 12437 11503 12495 11509
rect 12710 11500 12716 11552
rect 12768 11540 12774 11552
rect 12805 11543 12863 11549
rect 12805 11540 12817 11543
rect 12768 11512 12817 11540
rect 12768 11500 12774 11512
rect 12805 11509 12817 11512
rect 12851 11540 12863 11543
rect 13446 11540 13452 11552
rect 12851 11512 13452 11540
rect 12851 11509 12863 11512
rect 12805 11503 12863 11509
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 16482 11500 16488 11552
rect 16540 11540 16546 11552
rect 16853 11543 16911 11549
rect 16853 11540 16865 11543
rect 16540 11512 16865 11540
rect 16540 11500 16546 11512
rect 16853 11509 16865 11512
rect 16899 11509 16911 11543
rect 16853 11503 16911 11509
rect 18230 11500 18236 11552
rect 18288 11540 18294 11552
rect 18506 11540 18512 11552
rect 18288 11512 18512 11540
rect 18288 11500 18294 11512
rect 18506 11500 18512 11512
rect 18564 11500 18570 11552
rect 19306 11540 19334 11580
rect 19426 11568 19432 11620
rect 19484 11608 19490 11620
rect 19613 11611 19671 11617
rect 19613 11608 19625 11611
rect 19484 11580 19625 11608
rect 19484 11568 19490 11580
rect 19613 11577 19625 11580
rect 19659 11608 19671 11611
rect 19702 11608 19708 11620
rect 19659 11580 19708 11608
rect 19659 11577 19671 11580
rect 19613 11571 19671 11577
rect 19702 11568 19708 11580
rect 19760 11568 19766 11620
rect 19889 11611 19947 11617
rect 19889 11577 19901 11611
rect 19935 11608 19947 11611
rect 19978 11608 19984 11620
rect 19935 11580 19984 11608
rect 19935 11577 19947 11580
rect 19889 11571 19947 11577
rect 19904 11540 19932 11571
rect 19978 11568 19984 11580
rect 20036 11608 20042 11620
rect 21450 11608 21456 11620
rect 20036 11580 21456 11608
rect 20036 11568 20042 11580
rect 21450 11568 21456 11580
rect 21508 11568 21514 11620
rect 31389 11611 31447 11617
rect 31389 11577 31401 11611
rect 31435 11608 31447 11611
rect 31726 11608 31754 11648
rect 32582 11636 32588 11688
rect 32640 11676 32646 11688
rect 32677 11679 32735 11685
rect 32677 11676 32689 11679
rect 32640 11648 32689 11676
rect 32640 11636 32646 11648
rect 32677 11645 32689 11648
rect 32723 11645 32735 11679
rect 32677 11639 32735 11645
rect 31435 11580 31754 11608
rect 31435 11577 31447 11580
rect 31389 11571 31447 11577
rect 25682 11540 25688 11552
rect 19306 11512 19932 11540
rect 25643 11512 25688 11540
rect 25682 11500 25688 11512
rect 25740 11500 25746 11552
rect 26973 11543 27031 11549
rect 26973 11509 26985 11543
rect 27019 11540 27031 11543
rect 27338 11540 27344 11552
rect 27019 11512 27344 11540
rect 27019 11509 27031 11512
rect 26973 11503 27031 11509
rect 27338 11500 27344 11512
rect 27396 11500 27402 11552
rect 33318 11500 33324 11552
rect 33376 11540 33382 11552
rect 34517 11543 34575 11549
rect 34517 11540 34529 11543
rect 33376 11512 34529 11540
rect 33376 11500 33382 11512
rect 34517 11509 34529 11512
rect 34563 11509 34575 11543
rect 34517 11503 34575 11509
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 15565 11339 15623 11345
rect 15565 11305 15577 11339
rect 15611 11336 15623 11339
rect 15838 11336 15844 11348
rect 15611 11308 15844 11336
rect 15611 11305 15623 11308
rect 15565 11299 15623 11305
rect 15838 11296 15844 11308
rect 15896 11296 15902 11348
rect 18049 11339 18107 11345
rect 18049 11336 18061 11339
rect 16960 11308 18061 11336
rect 13446 11268 13452 11280
rect 13359 11240 13452 11268
rect 13446 11228 13452 11240
rect 13504 11268 13510 11280
rect 16393 11271 16451 11277
rect 13504 11240 15700 11268
rect 13504 11228 13510 11240
rect 15672 11212 15700 11240
rect 16393 11237 16405 11271
rect 16439 11268 16451 11271
rect 16850 11268 16856 11280
rect 16439 11240 16856 11268
rect 16439 11237 16451 11240
rect 16393 11231 16451 11237
rect 16850 11228 16856 11240
rect 16908 11228 16914 11280
rect 14737 11203 14795 11209
rect 14737 11169 14749 11203
rect 14783 11200 14795 11203
rect 15562 11200 15568 11212
rect 14783 11172 15568 11200
rect 14783 11169 14795 11172
rect 14737 11163 14795 11169
rect 15562 11160 15568 11172
rect 15620 11160 15626 11212
rect 15654 11160 15660 11212
rect 15712 11200 15718 11212
rect 16960 11209 16988 11308
rect 18049 11305 18061 11308
rect 18095 11305 18107 11339
rect 18049 11299 18107 11305
rect 18322 11296 18328 11348
rect 18380 11336 18386 11348
rect 18417 11339 18475 11345
rect 18417 11336 18429 11339
rect 18380 11308 18429 11336
rect 18380 11296 18386 11308
rect 18417 11305 18429 11308
rect 18463 11305 18475 11339
rect 18417 11299 18475 11305
rect 20254 11296 20260 11348
rect 20312 11336 20318 11348
rect 20625 11339 20683 11345
rect 20625 11336 20637 11339
rect 20312 11308 20637 11336
rect 20312 11296 20318 11308
rect 20625 11305 20637 11308
rect 20671 11305 20683 11339
rect 20625 11299 20683 11305
rect 21082 11296 21088 11348
rect 21140 11336 21146 11348
rect 21361 11339 21419 11345
rect 21361 11336 21373 11339
rect 21140 11308 21373 11336
rect 21140 11296 21146 11308
rect 21361 11305 21373 11308
rect 21407 11305 21419 11339
rect 21361 11299 21419 11305
rect 21450 11296 21456 11348
rect 21508 11336 21514 11348
rect 23014 11336 23020 11348
rect 21508 11308 23020 11336
rect 21508 11296 21514 11308
rect 23014 11296 23020 11308
rect 23072 11296 23078 11348
rect 25498 11296 25504 11348
rect 25556 11336 25562 11348
rect 25777 11339 25835 11345
rect 25777 11336 25789 11339
rect 25556 11308 25789 11336
rect 25556 11296 25562 11308
rect 25777 11305 25789 11308
rect 25823 11305 25835 11339
rect 25777 11299 25835 11305
rect 27890 11296 27896 11348
rect 27948 11336 27954 11348
rect 28537 11339 28595 11345
rect 28537 11336 28549 11339
rect 27948 11308 28549 11336
rect 27948 11296 27954 11308
rect 28537 11305 28549 11308
rect 28583 11305 28595 11339
rect 28537 11299 28595 11305
rect 30024 11308 31754 11336
rect 17221 11271 17279 11277
rect 17221 11237 17233 11271
rect 17267 11237 17279 11271
rect 17221 11231 17279 11237
rect 17405 11271 17463 11277
rect 17405 11237 17417 11271
rect 17451 11268 17463 11271
rect 18230 11268 18236 11280
rect 17451 11240 18236 11268
rect 17451 11237 17463 11240
rect 17405 11231 17463 11237
rect 16945 11203 17003 11209
rect 16945 11200 16957 11203
rect 15712 11172 16957 11200
rect 15712 11160 15718 11172
rect 16945 11169 16957 11172
rect 16991 11169 17003 11203
rect 16945 11163 17003 11169
rect 9953 11135 10011 11141
rect 9953 11101 9965 11135
rect 9999 11101 10011 11135
rect 9953 11095 10011 11101
rect 10137 11135 10195 11141
rect 10137 11101 10149 11135
rect 10183 11132 10195 11135
rect 10410 11132 10416 11144
rect 10183 11104 10416 11132
rect 10183 11101 10195 11104
rect 10137 11095 10195 11101
rect 9968 11064 9996 11095
rect 10410 11092 10416 11104
rect 10468 11092 10474 11144
rect 11514 11092 11520 11144
rect 11572 11132 11578 11144
rect 12342 11141 12348 11144
rect 12069 11135 12127 11141
rect 12069 11132 12081 11135
rect 11572 11104 12081 11132
rect 11572 11092 11578 11104
rect 12069 11101 12081 11104
rect 12115 11101 12127 11135
rect 12336 11132 12348 11141
rect 12303 11104 12348 11132
rect 12069 11095 12127 11101
rect 12336 11095 12348 11104
rect 12342 11092 12348 11095
rect 12400 11092 12406 11144
rect 14274 11092 14280 11144
rect 14332 11132 14338 11144
rect 14553 11135 14611 11141
rect 14553 11132 14565 11135
rect 14332 11104 14565 11132
rect 14332 11092 14338 11104
rect 14553 11101 14565 11104
rect 14599 11101 14611 11135
rect 14553 11095 14611 11101
rect 15286 11092 15292 11144
rect 15344 11132 15350 11144
rect 17236 11132 17264 11231
rect 18230 11228 18236 11240
rect 18288 11228 18294 11280
rect 21910 11228 21916 11280
rect 21968 11268 21974 11280
rect 21968 11240 23336 11268
rect 21968 11228 21974 11240
rect 18138 11160 18144 11212
rect 18196 11200 18202 11212
rect 18598 11200 18604 11212
rect 18196 11172 18604 11200
rect 18196 11160 18202 11172
rect 18598 11160 18604 11172
rect 18656 11160 18662 11212
rect 23308 11209 23336 11240
rect 23474 11228 23480 11280
rect 23532 11268 23538 11280
rect 24394 11268 24400 11280
rect 23532 11240 24400 11268
rect 23532 11228 23538 11240
rect 24394 11228 24400 11240
rect 24452 11228 24458 11280
rect 23293 11203 23351 11209
rect 23293 11169 23305 11203
rect 23339 11200 23351 11203
rect 24118 11200 24124 11212
rect 23339 11172 24124 11200
rect 23339 11169 23351 11172
rect 23293 11163 23351 11169
rect 24118 11160 24124 11172
rect 24176 11160 24182 11212
rect 29914 11160 29920 11212
rect 29972 11200 29978 11212
rect 30024 11209 30052 11308
rect 31726 11268 31754 11308
rect 32582 11268 32588 11280
rect 31726 11240 32588 11268
rect 32582 11228 32588 11240
rect 32640 11268 32646 11280
rect 33689 11271 33747 11277
rect 33689 11268 33701 11271
rect 32640 11240 33701 11268
rect 32640 11228 32646 11240
rect 33689 11237 33701 11240
rect 33735 11237 33747 11271
rect 33689 11231 33747 11237
rect 30009 11203 30067 11209
rect 30009 11200 30021 11203
rect 29972 11172 30021 11200
rect 29972 11160 29978 11172
rect 30009 11169 30021 11172
rect 30055 11169 30067 11203
rect 30009 11163 30067 11169
rect 17957 11135 18015 11141
rect 17957 11132 17969 11135
rect 15344 11104 17969 11132
rect 15344 11092 15350 11104
rect 17957 11101 17969 11104
rect 18003 11101 18015 11135
rect 19242 11132 19248 11144
rect 19203 11104 19248 11132
rect 17957 11095 18015 11101
rect 19242 11092 19248 11104
rect 19300 11092 19306 11144
rect 19794 11092 19800 11144
rect 19852 11132 19858 11144
rect 21082 11132 21088 11144
rect 19852 11104 21088 11132
rect 19852 11092 19858 11104
rect 21082 11092 21088 11104
rect 21140 11132 21146 11144
rect 21358 11141 21364 11144
rect 21177 11135 21235 11141
rect 21177 11132 21189 11135
rect 21140 11104 21189 11132
rect 21140 11092 21146 11104
rect 21177 11101 21189 11104
rect 21223 11101 21235 11135
rect 21177 11095 21235 11101
rect 21315 11135 21364 11141
rect 21315 11101 21327 11135
rect 21361 11101 21364 11135
rect 21315 11095 21364 11101
rect 21358 11092 21364 11095
rect 21416 11092 21422 11144
rect 21545 11135 21603 11141
rect 21545 11132 21557 11135
rect 21468 11104 21557 11132
rect 10778 11064 10784 11076
rect 9968 11036 10784 11064
rect 10778 11024 10784 11036
rect 10836 11024 10842 11076
rect 13814 11024 13820 11076
rect 13872 11064 13878 11076
rect 14369 11067 14427 11073
rect 14369 11064 14381 11067
rect 13872 11036 14381 11064
rect 13872 11024 13878 11036
rect 14369 11033 14381 11036
rect 14415 11033 14427 11067
rect 15194 11064 15200 11076
rect 15155 11036 15200 11064
rect 14369 11027 14427 11033
rect 15194 11024 15200 11036
rect 15252 11024 15258 11076
rect 15381 11067 15439 11073
rect 15381 11033 15393 11067
rect 15427 11064 15439 11067
rect 15562 11064 15568 11076
rect 15427 11036 15568 11064
rect 15427 11033 15439 11036
rect 15381 11027 15439 11033
rect 15562 11024 15568 11036
rect 15620 11064 15626 11076
rect 15620 11036 15976 11064
rect 15620 11024 15626 11036
rect 10042 10996 10048 11008
rect 10003 10968 10048 10996
rect 10042 10956 10048 10968
rect 10100 10956 10106 11008
rect 15948 10996 15976 11036
rect 16022 11024 16028 11076
rect 16080 11064 16086 11076
rect 16209 11067 16267 11073
rect 16080 11036 16125 11064
rect 16080 11024 16086 11036
rect 16209 11033 16221 11067
rect 16255 11033 16267 11067
rect 16209 11027 16267 11033
rect 19512 11067 19570 11073
rect 19512 11033 19524 11067
rect 19558 11064 19570 11067
rect 20070 11064 20076 11076
rect 19558 11036 20076 11064
rect 19558 11033 19570 11036
rect 19512 11027 19570 11033
rect 16224 10996 16252 11027
rect 20070 11024 20076 11036
rect 20128 11024 20134 11076
rect 20530 11024 20536 11076
rect 20588 11064 20594 11076
rect 20588 11036 21312 11064
rect 20588 11024 20594 11036
rect 15948 10968 16252 10996
rect 19334 10956 19340 11008
rect 19392 10996 19398 11008
rect 20254 10996 20260 11008
rect 19392 10968 20260 10996
rect 19392 10956 19398 10968
rect 20254 10956 20260 10968
rect 20312 10956 20318 11008
rect 21284 10996 21312 11036
rect 21468 10996 21496 11104
rect 21545 11101 21557 11104
rect 21591 11101 21603 11135
rect 23014 11132 23020 11144
rect 22975 11104 23020 11132
rect 21545 11095 21603 11101
rect 23014 11092 23020 11104
rect 23072 11092 23078 11144
rect 24397 11135 24455 11141
rect 24397 11101 24409 11135
rect 24443 11132 24455 11135
rect 25590 11132 25596 11144
rect 24443 11104 25596 11132
rect 24443 11101 24455 11104
rect 24397 11095 24455 11101
rect 25590 11092 25596 11104
rect 25648 11092 25654 11144
rect 26234 11092 26240 11144
rect 26292 11132 26298 11144
rect 27157 11135 27215 11141
rect 27157 11132 27169 11135
rect 26292 11104 27169 11132
rect 26292 11092 26298 11104
rect 27157 11101 27169 11104
rect 27203 11101 27215 11135
rect 32398 11132 32404 11144
rect 32311 11104 32404 11132
rect 27157 11095 27215 11101
rect 32398 11092 32404 11104
rect 32456 11132 32462 11144
rect 34698 11132 34704 11144
rect 32456 11104 34704 11132
rect 32456 11092 32462 11104
rect 34698 11092 34704 11104
rect 34756 11092 34762 11144
rect 24664 11067 24722 11073
rect 24664 11033 24676 11067
rect 24710 11064 24722 11067
rect 25682 11064 25688 11076
rect 24710 11036 25688 11064
rect 24710 11033 24722 11036
rect 24664 11027 24722 11033
rect 25682 11024 25688 11036
rect 25740 11024 25746 11076
rect 27424 11067 27482 11073
rect 27424 11033 27436 11067
rect 27470 11064 27482 11067
rect 27522 11064 27528 11076
rect 27470 11036 27528 11064
rect 27470 11033 27482 11036
rect 27424 11027 27482 11033
rect 27522 11024 27528 11036
rect 27580 11024 27586 11076
rect 30276 11067 30334 11073
rect 30276 11033 30288 11067
rect 30322 11064 30334 11067
rect 30926 11064 30932 11076
rect 30322 11036 30932 11064
rect 30322 11033 30334 11036
rect 30276 11027 30334 11033
rect 30926 11024 30932 11036
rect 30984 11024 30990 11076
rect 21284 10968 21496 10996
rect 30374 10956 30380 11008
rect 30432 10996 30438 11008
rect 30834 10996 30840 11008
rect 30432 10968 30840 10996
rect 30432 10956 30438 10968
rect 30834 10956 30840 10968
rect 30892 10996 30898 11008
rect 31389 10999 31447 11005
rect 31389 10996 31401 10999
rect 30892 10968 31401 10996
rect 30892 10956 30898 10968
rect 31389 10965 31401 10968
rect 31435 10965 31447 10999
rect 31389 10959 31447 10965
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 7558 10752 7564 10804
rect 7616 10792 7622 10804
rect 10318 10792 10324 10804
rect 7616 10764 10324 10792
rect 7616 10752 7622 10764
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 14553 10795 14611 10801
rect 14553 10761 14565 10795
rect 14599 10792 14611 10795
rect 16390 10792 16396 10804
rect 14599 10764 16396 10792
rect 14599 10761 14611 10764
rect 14553 10755 14611 10761
rect 16390 10752 16396 10764
rect 16448 10752 16454 10804
rect 16666 10752 16672 10804
rect 16724 10792 16730 10804
rect 17129 10795 17187 10801
rect 17129 10792 17141 10795
rect 16724 10764 17141 10792
rect 16724 10752 16730 10764
rect 17129 10761 17141 10764
rect 17175 10761 17187 10795
rect 17129 10755 17187 10761
rect 17218 10752 17224 10804
rect 17276 10792 17282 10804
rect 20070 10792 20076 10804
rect 17276 10764 19564 10792
rect 20031 10764 20076 10792
rect 17276 10752 17282 10764
rect 8680 10696 11100 10724
rect 8680 10665 8708 10696
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 8932 10659 8990 10665
rect 8932 10625 8944 10659
rect 8978 10656 8990 10659
rect 10042 10656 10048 10668
rect 8978 10628 10048 10656
rect 8978 10625 8990 10628
rect 8932 10619 8990 10625
rect 10042 10616 10048 10628
rect 10100 10616 10106 10668
rect 10318 10616 10324 10668
rect 10376 10656 10382 10668
rect 10965 10659 11023 10665
rect 10965 10656 10977 10659
rect 10376 10628 10977 10656
rect 10376 10616 10382 10628
rect 10965 10625 10977 10628
rect 11011 10625 11023 10659
rect 11072 10656 11100 10696
rect 15010 10684 15016 10736
rect 15068 10724 15074 10736
rect 16117 10727 16175 10733
rect 16117 10724 16129 10727
rect 15068 10696 16129 10724
rect 15068 10684 15074 10696
rect 16117 10693 16129 10696
rect 16163 10693 16175 10727
rect 18874 10724 18880 10736
rect 16117 10687 16175 10693
rect 16776 10696 18880 10724
rect 16776 10668 16804 10696
rect 18874 10684 18880 10696
rect 18932 10684 18938 10736
rect 19153 10727 19211 10733
rect 19153 10693 19165 10727
rect 19199 10724 19211 10727
rect 19426 10724 19432 10736
rect 19199 10696 19432 10724
rect 19199 10693 19211 10696
rect 19153 10687 19211 10693
rect 19426 10684 19432 10696
rect 19484 10684 19490 10736
rect 19536 10724 19564 10764
rect 20070 10752 20076 10764
rect 20128 10752 20134 10804
rect 21082 10752 21088 10804
rect 21140 10792 21146 10804
rect 27614 10792 27620 10804
rect 21140 10764 22784 10792
rect 21140 10752 21146 10764
rect 22756 10736 22784 10764
rect 25148 10764 27620 10792
rect 19536 10696 22094 10724
rect 11514 10656 11520 10668
rect 11072 10628 11520 10656
rect 10965 10619 11023 10625
rect 11514 10616 11520 10628
rect 11572 10616 11578 10668
rect 11606 10616 11612 10668
rect 11664 10656 11670 10668
rect 11773 10659 11831 10665
rect 11773 10656 11785 10659
rect 11664 10628 11785 10656
rect 11664 10616 11670 10628
rect 11773 10625 11785 10628
rect 11819 10625 11831 10659
rect 13998 10656 14004 10668
rect 13959 10628 14004 10656
rect 11773 10619 11831 10625
rect 13998 10616 14004 10628
rect 14056 10616 14062 10668
rect 15105 10659 15163 10665
rect 15105 10625 15117 10659
rect 15151 10656 15163 10659
rect 15286 10656 15292 10668
rect 15151 10628 15292 10656
rect 15151 10625 15163 10628
rect 15105 10619 15163 10625
rect 10781 10591 10839 10597
rect 10781 10588 10793 10591
rect 10060 10560 10793 10588
rect 10060 10529 10088 10560
rect 10781 10557 10793 10560
rect 10827 10588 10839 10591
rect 11422 10588 11428 10600
rect 10827 10560 11428 10588
rect 10827 10557 10839 10560
rect 10781 10551 10839 10557
rect 11422 10548 11428 10560
rect 11480 10548 11486 10600
rect 14274 10588 14280 10600
rect 14235 10560 14280 10588
rect 14274 10548 14280 10560
rect 14332 10548 14338 10600
rect 10045 10523 10103 10529
rect 10045 10489 10057 10523
rect 10091 10489 10103 10523
rect 10594 10520 10600 10532
rect 10555 10492 10600 10520
rect 10045 10483 10103 10489
rect 10594 10480 10600 10492
rect 10652 10480 10658 10532
rect 10870 10520 10876 10532
rect 10831 10492 10876 10520
rect 10870 10480 10876 10492
rect 10928 10480 10934 10532
rect 12894 10520 12900 10532
rect 12807 10492 12900 10520
rect 12894 10480 12900 10492
rect 12952 10520 12958 10532
rect 15120 10520 15148 10619
rect 15286 10616 15292 10628
rect 15344 10616 15350 10668
rect 15565 10659 15623 10665
rect 15565 10625 15577 10659
rect 15611 10656 15623 10659
rect 15654 10656 15660 10668
rect 15611 10628 15660 10656
rect 15611 10625 15623 10628
rect 15565 10619 15623 10625
rect 15654 10616 15660 10628
rect 15712 10616 15718 10668
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10656 15991 10659
rect 16206 10656 16212 10668
rect 15979 10628 16212 10656
rect 15979 10625 15991 10628
rect 15933 10619 15991 10625
rect 16206 10616 16212 10628
rect 16264 10616 16270 10668
rect 16669 10659 16727 10665
rect 16669 10625 16681 10659
rect 16715 10625 16727 10659
rect 16669 10619 16727 10625
rect 15194 10548 15200 10600
rect 15252 10588 15258 10600
rect 16684 10588 16712 10619
rect 16758 10616 16764 10668
rect 16816 10656 16822 10668
rect 16945 10659 17003 10665
rect 16816 10628 16909 10656
rect 16816 10616 16822 10628
rect 16945 10625 16957 10659
rect 16991 10625 17003 10659
rect 16945 10619 17003 10625
rect 15252 10560 16712 10588
rect 15252 10548 15258 10560
rect 12952 10492 15148 10520
rect 12952 10480 12958 10492
rect 10778 10452 10784 10464
rect 10739 10424 10784 10452
rect 10778 10412 10784 10424
rect 10836 10412 10842 10464
rect 13814 10412 13820 10464
rect 13872 10452 13878 10464
rect 14093 10455 14151 10461
rect 14093 10452 14105 10455
rect 13872 10424 14105 10452
rect 13872 10412 13878 10424
rect 14093 10421 14105 10424
rect 14139 10421 14151 10455
rect 14093 10415 14151 10421
rect 16390 10412 16396 10464
rect 16448 10452 16454 10464
rect 16960 10452 16988 10619
rect 17586 10616 17592 10668
rect 17644 10656 17650 10668
rect 19521 10659 19579 10665
rect 19521 10656 19533 10659
rect 17644 10628 19533 10656
rect 17644 10616 17650 10628
rect 19521 10625 19533 10628
rect 19567 10625 19579 10659
rect 19521 10619 19579 10625
rect 19981 10659 20039 10665
rect 19981 10625 19993 10659
rect 20027 10625 20039 10659
rect 19981 10619 20039 10625
rect 20165 10659 20223 10665
rect 20165 10625 20177 10659
rect 20211 10656 20223 10659
rect 21266 10656 21272 10668
rect 20211 10628 21272 10656
rect 20211 10625 20223 10628
rect 20165 10619 20223 10625
rect 19334 10548 19340 10600
rect 19392 10588 19398 10600
rect 19392 10560 19437 10588
rect 19392 10548 19398 10560
rect 19996 10520 20024 10619
rect 21266 10616 21272 10628
rect 21324 10656 21330 10668
rect 21910 10656 21916 10668
rect 21324 10628 21916 10656
rect 21324 10616 21330 10628
rect 21910 10616 21916 10628
rect 21968 10616 21974 10668
rect 22066 10656 22094 10696
rect 22738 10684 22744 10736
rect 22796 10724 22802 10736
rect 24213 10727 24271 10733
rect 24213 10724 24225 10727
rect 22796 10696 24225 10724
rect 22796 10684 22802 10696
rect 24213 10693 24225 10696
rect 24259 10724 24271 10727
rect 24765 10727 24823 10733
rect 24765 10724 24777 10727
rect 24259 10696 24777 10724
rect 24259 10693 24271 10696
rect 24213 10687 24271 10693
rect 24765 10693 24777 10696
rect 24811 10693 24823 10727
rect 24765 10687 24823 10693
rect 25148 10665 25176 10764
rect 27614 10752 27620 10764
rect 27672 10752 27678 10804
rect 31018 10792 31024 10804
rect 27908 10764 31024 10792
rect 27798 10684 27804 10736
rect 27856 10684 27862 10736
rect 24029 10659 24087 10665
rect 24029 10656 24041 10659
rect 22066 10628 24041 10656
rect 24029 10625 24041 10628
rect 24075 10625 24087 10659
rect 24029 10619 24087 10625
rect 25133 10659 25191 10665
rect 25133 10625 25145 10659
rect 25179 10625 25191 10659
rect 25133 10619 25191 10625
rect 19352 10492 20024 10520
rect 24044 10520 24072 10619
rect 25314 10616 25320 10668
rect 25372 10656 25378 10668
rect 27663 10659 27721 10665
rect 25372 10628 27568 10656
rect 25372 10616 25378 10628
rect 24949 10591 25007 10597
rect 24949 10557 24961 10591
rect 24995 10588 25007 10591
rect 25498 10588 25504 10600
rect 24995 10560 25504 10588
rect 24995 10557 25007 10560
rect 24949 10551 25007 10557
rect 25498 10548 25504 10560
rect 25556 10548 25562 10600
rect 27540 10588 27568 10628
rect 27663 10625 27675 10659
rect 27709 10656 27721 10659
rect 27816 10656 27844 10684
rect 27908 10665 27936 10764
rect 31018 10752 31024 10764
rect 31076 10752 31082 10804
rect 33226 10752 33232 10804
rect 33284 10792 33290 10804
rect 34057 10795 34115 10801
rect 34057 10792 34069 10795
rect 33284 10764 34069 10792
rect 33284 10752 33290 10764
rect 34057 10761 34069 10764
rect 34103 10761 34115 10795
rect 34057 10755 34115 10761
rect 29546 10724 29552 10736
rect 28966 10696 29552 10724
rect 27709 10628 27844 10656
rect 27893 10659 27951 10665
rect 27709 10625 27721 10628
rect 27663 10619 27721 10625
rect 27893 10625 27905 10659
rect 27939 10625 27951 10659
rect 27893 10619 27951 10625
rect 27801 10591 27859 10597
rect 27801 10588 27813 10591
rect 27540 10560 27813 10588
rect 27801 10557 27813 10560
rect 27847 10588 27859 10591
rect 28966 10588 28994 10696
rect 29546 10684 29552 10696
rect 29604 10684 29610 10736
rect 30466 10684 30472 10736
rect 30524 10724 30530 10736
rect 30723 10727 30781 10733
rect 30723 10724 30735 10727
rect 30524 10696 30735 10724
rect 30524 10684 30530 10696
rect 30723 10693 30735 10696
rect 30769 10693 30781 10727
rect 32766 10724 32772 10736
rect 30723 10687 30781 10693
rect 31726 10696 32772 10724
rect 29362 10616 29368 10668
rect 29420 10665 29426 10668
rect 29420 10659 29469 10665
rect 29420 10625 29423 10659
rect 29457 10625 29469 10659
rect 29420 10619 29469 10625
rect 29641 10659 29699 10665
rect 29641 10625 29653 10659
rect 29687 10656 29699 10659
rect 30558 10656 30564 10668
rect 29687 10628 30564 10656
rect 29687 10625 29699 10628
rect 29641 10619 29699 10625
rect 29420 10616 29426 10619
rect 30558 10616 30564 10628
rect 30616 10616 30622 10668
rect 31021 10659 31079 10665
rect 31021 10625 31033 10659
rect 31067 10656 31079 10659
rect 31726 10656 31754 10696
rect 32766 10684 32772 10696
rect 32824 10684 32830 10736
rect 32944 10727 33002 10733
rect 32944 10693 32956 10727
rect 32990 10724 33002 10727
rect 33318 10724 33324 10736
rect 32990 10696 33324 10724
rect 32990 10693 33002 10696
rect 32944 10687 33002 10693
rect 33318 10684 33324 10696
rect 33376 10684 33382 10736
rect 31067 10628 31754 10656
rect 31067 10625 31079 10628
rect 31021 10619 31079 10625
rect 30834 10588 30840 10600
rect 27847 10560 28994 10588
rect 30795 10560 30840 10588
rect 27847 10557 27859 10560
rect 27801 10551 27859 10557
rect 30834 10548 30840 10560
rect 30892 10548 30898 10600
rect 32582 10548 32588 10600
rect 32640 10588 32646 10600
rect 32677 10591 32735 10597
rect 32677 10588 32689 10591
rect 32640 10560 32689 10588
rect 32640 10548 32646 10560
rect 32677 10557 32689 10560
rect 32723 10557 32735 10591
rect 32677 10551 32735 10557
rect 24044 10492 25636 10520
rect 19352 10461 19380 10492
rect 25608 10464 25636 10492
rect 26970 10480 26976 10532
rect 27028 10520 27034 10532
rect 27525 10523 27583 10529
rect 27525 10520 27537 10523
rect 27028 10492 27537 10520
rect 27028 10480 27034 10492
rect 27525 10489 27537 10492
rect 27571 10520 27583 10523
rect 29273 10523 29331 10529
rect 29273 10520 29285 10523
rect 27571 10492 29285 10520
rect 27571 10489 27583 10492
rect 27525 10483 27583 10489
rect 29273 10489 29285 10492
rect 29319 10520 29331 10523
rect 30374 10520 30380 10532
rect 29319 10492 30380 10520
rect 29319 10489 29331 10492
rect 29273 10483 29331 10489
rect 30374 10480 30380 10492
rect 30432 10520 30438 10532
rect 30653 10523 30711 10529
rect 30653 10520 30665 10523
rect 30432 10492 30665 10520
rect 30432 10480 30438 10492
rect 30653 10489 30665 10492
rect 30699 10489 30711 10523
rect 30653 10483 30711 10489
rect 16448 10424 16988 10452
rect 19337 10455 19395 10461
rect 16448 10412 16454 10424
rect 19337 10421 19349 10455
rect 19383 10421 19395 10455
rect 19337 10415 19395 10421
rect 19429 10455 19487 10461
rect 19429 10421 19441 10455
rect 19475 10452 19487 10455
rect 19978 10452 19984 10464
rect 19475 10424 19984 10452
rect 19475 10421 19487 10424
rect 19429 10415 19487 10421
rect 19978 10412 19984 10424
rect 20036 10412 20042 10464
rect 24946 10452 24952 10464
rect 24907 10424 24952 10452
rect 24946 10412 24952 10424
rect 25004 10412 25010 10464
rect 25041 10455 25099 10461
rect 25041 10421 25053 10455
rect 25087 10452 25099 10455
rect 25314 10452 25320 10464
rect 25087 10424 25320 10452
rect 25087 10421 25099 10424
rect 25041 10415 25099 10421
rect 25314 10412 25320 10424
rect 25372 10412 25378 10464
rect 25590 10412 25596 10464
rect 25648 10452 25654 10464
rect 26694 10452 26700 10464
rect 25648 10424 26700 10452
rect 25648 10412 25654 10424
rect 26694 10412 26700 10424
rect 26752 10412 26758 10464
rect 27430 10412 27436 10464
rect 27488 10452 27494 10464
rect 27709 10455 27767 10461
rect 27709 10452 27721 10455
rect 27488 10424 27721 10452
rect 27488 10412 27494 10424
rect 27709 10421 27721 10424
rect 27755 10421 27767 10455
rect 27709 10415 27767 10421
rect 28810 10412 28816 10464
rect 28868 10452 28874 10464
rect 29457 10455 29515 10461
rect 29457 10452 29469 10455
rect 28868 10424 29469 10452
rect 28868 10412 28874 10424
rect 29457 10421 29469 10424
rect 29503 10421 29515 10455
rect 29457 10415 29515 10421
rect 29546 10412 29552 10464
rect 29604 10452 29610 10464
rect 30929 10455 30987 10461
rect 30929 10452 30941 10455
rect 29604 10424 30941 10452
rect 29604 10412 29610 10424
rect 30929 10421 30941 10424
rect 30975 10452 30987 10455
rect 31110 10452 31116 10464
rect 30975 10424 31116 10452
rect 30975 10421 30987 10424
rect 30929 10415 30987 10421
rect 31110 10412 31116 10424
rect 31168 10412 31174 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 10965 10251 11023 10257
rect 10965 10217 10977 10251
rect 11011 10248 11023 10251
rect 11606 10248 11612 10260
rect 11011 10220 11612 10248
rect 11011 10217 11023 10220
rect 10965 10211 11023 10217
rect 11606 10208 11612 10220
rect 11664 10208 11670 10260
rect 14274 10208 14280 10260
rect 14332 10248 14338 10260
rect 14645 10251 14703 10257
rect 14645 10248 14657 10251
rect 14332 10220 14657 10248
rect 14332 10208 14338 10220
rect 14645 10217 14657 10220
rect 14691 10217 14703 10251
rect 14645 10211 14703 10217
rect 15013 10251 15071 10257
rect 15013 10217 15025 10251
rect 15059 10248 15071 10251
rect 15194 10248 15200 10260
rect 15059 10220 15200 10248
rect 15059 10217 15071 10220
rect 15013 10211 15071 10217
rect 15194 10208 15200 10220
rect 15252 10208 15258 10260
rect 16482 10248 16488 10260
rect 16443 10220 16488 10248
rect 16482 10208 16488 10220
rect 16540 10208 16546 10260
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 18601 10251 18659 10257
rect 18601 10248 18613 10251
rect 18012 10220 18613 10248
rect 18012 10208 18018 10220
rect 18601 10217 18613 10220
rect 18647 10248 18659 10251
rect 18690 10248 18696 10260
rect 18647 10220 18696 10248
rect 18647 10217 18659 10220
rect 18601 10211 18659 10217
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 25866 10208 25872 10260
rect 25924 10248 25930 10260
rect 26973 10251 27031 10257
rect 26973 10248 26985 10251
rect 25924 10220 26985 10248
rect 25924 10208 25930 10220
rect 26973 10217 26985 10220
rect 27019 10217 27031 10251
rect 27522 10248 27528 10260
rect 27483 10220 27528 10248
rect 26973 10211 27031 10217
rect 27522 10208 27528 10220
rect 27580 10208 27586 10260
rect 30926 10248 30932 10260
rect 30887 10220 30932 10248
rect 30926 10208 30932 10220
rect 30984 10208 30990 10260
rect 33594 10208 33600 10260
rect 33652 10248 33658 10260
rect 34057 10251 34115 10257
rect 34057 10248 34069 10251
rect 33652 10220 34069 10248
rect 33652 10208 33658 10220
rect 34057 10217 34069 10220
rect 34103 10217 34115 10251
rect 34057 10211 34115 10217
rect 10594 10140 10600 10192
rect 10652 10180 10658 10192
rect 14090 10180 14096 10192
rect 10652 10152 14096 10180
rect 10652 10140 10658 10152
rect 14090 10140 14096 10152
rect 14148 10180 14154 10192
rect 15749 10183 15807 10189
rect 15749 10180 15761 10183
rect 14148 10152 15761 10180
rect 14148 10140 14154 10152
rect 15749 10149 15761 10152
rect 15795 10149 15807 10183
rect 15749 10143 15807 10149
rect 17218 10140 17224 10192
rect 17276 10140 17282 10192
rect 26694 10140 26700 10192
rect 26752 10180 26758 10192
rect 32674 10180 32680 10192
rect 26752 10152 32680 10180
rect 26752 10140 26758 10152
rect 10686 10072 10692 10124
rect 10744 10112 10750 10124
rect 10781 10115 10839 10121
rect 10781 10112 10793 10115
rect 10744 10084 10793 10112
rect 10744 10072 10750 10084
rect 10781 10081 10793 10084
rect 10827 10081 10839 10115
rect 12894 10112 12900 10124
rect 10781 10075 10839 10081
rect 12820 10084 12900 10112
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10044 1915 10047
rect 9122 10044 9128 10056
rect 1903 10016 2774 10044
rect 9083 10016 9128 10044
rect 1903 10013 1915 10016
rect 1857 10007 1915 10013
rect 2746 9976 2774 10016
rect 9122 10004 9128 10016
rect 9180 10004 9186 10056
rect 10870 10004 10876 10056
rect 10928 10044 10934 10056
rect 11241 10047 11299 10053
rect 11241 10044 11253 10047
rect 10928 10016 11253 10044
rect 10928 10004 10934 10016
rect 11241 10013 11253 10016
rect 11287 10013 11299 10047
rect 11241 10007 11299 10013
rect 11330 10004 11336 10056
rect 11388 10044 11394 10056
rect 12621 10047 12679 10053
rect 11388 10016 12434 10044
rect 11388 10004 11394 10016
rect 12406 9976 12434 10016
rect 12621 10013 12633 10047
rect 12667 10044 12679 10047
rect 12710 10044 12716 10056
rect 12667 10016 12716 10044
rect 12667 10013 12679 10016
rect 12621 10007 12679 10013
rect 12710 10004 12716 10016
rect 12768 10004 12774 10056
rect 12820 10053 12848 10084
rect 12894 10072 12900 10084
rect 12952 10072 12958 10124
rect 13998 10072 14004 10124
rect 14056 10112 14062 10124
rect 14737 10115 14795 10121
rect 14737 10112 14749 10115
rect 14056 10084 14749 10112
rect 14056 10072 14062 10084
rect 14737 10081 14749 10084
rect 14783 10081 14795 10115
rect 17236 10112 17264 10140
rect 29564 10121 29592 10152
rect 32674 10140 32680 10152
rect 32732 10140 32738 10192
rect 14737 10075 14795 10081
rect 15580 10084 17264 10112
rect 29549 10115 29607 10121
rect 12805 10047 12863 10053
rect 12805 10013 12817 10047
rect 12851 10013 12863 10047
rect 12805 10007 12863 10013
rect 13814 10004 13820 10056
rect 13872 10044 13878 10056
rect 15580 10053 15608 10084
rect 29549 10081 29561 10115
rect 29595 10081 29607 10115
rect 29549 10075 29607 10081
rect 29825 10115 29883 10121
rect 29825 10081 29837 10115
rect 29871 10112 29883 10115
rect 30374 10112 30380 10124
rect 29871 10084 30380 10112
rect 29871 10081 29883 10084
rect 29825 10075 29883 10081
rect 30374 10072 30380 10084
rect 30432 10072 30438 10124
rect 32232 10084 32812 10112
rect 14645 10047 14703 10053
rect 14645 10044 14657 10047
rect 13872 10016 14657 10044
rect 13872 10004 13878 10016
rect 14645 10013 14657 10016
rect 14691 10013 14703 10047
rect 14645 10007 14703 10013
rect 15565 10047 15623 10053
rect 15565 10013 15577 10047
rect 15611 10013 15623 10047
rect 15565 10007 15623 10013
rect 16114 10004 16120 10056
rect 16172 10044 16178 10056
rect 17221 10047 17279 10053
rect 17221 10044 17233 10047
rect 16172 10016 17233 10044
rect 16172 10004 16178 10016
rect 17221 10013 17233 10016
rect 17267 10013 17279 10047
rect 17221 10007 17279 10013
rect 19334 10004 19340 10056
rect 19392 10044 19398 10056
rect 20533 10047 20591 10053
rect 20533 10044 20545 10047
rect 19392 10016 20545 10044
rect 19392 10004 19398 10016
rect 20533 10013 20545 10016
rect 20579 10044 20591 10047
rect 21910 10044 21916 10056
rect 20579 10016 21916 10044
rect 20579 10013 20591 10016
rect 20533 10007 20591 10013
rect 21910 10004 21916 10016
rect 21968 10004 21974 10056
rect 23014 10004 23020 10056
rect 23072 10044 23078 10056
rect 24857 10047 24915 10053
rect 24857 10044 24869 10047
rect 23072 10016 24869 10044
rect 23072 10004 23078 10016
rect 24857 10013 24869 10016
rect 24903 10013 24915 10047
rect 24857 10007 24915 10013
rect 25593 10047 25651 10053
rect 25593 10013 25605 10047
rect 25639 10044 25651 10047
rect 26234 10044 26240 10056
rect 25639 10016 26240 10044
rect 25639 10013 25651 10016
rect 25593 10007 25651 10013
rect 26234 10004 26240 10016
rect 26292 10004 26298 10056
rect 27430 10044 27436 10056
rect 27391 10016 27436 10044
rect 27430 10004 27436 10016
rect 27488 10004 27494 10056
rect 27617 10047 27675 10053
rect 27617 10013 27629 10047
rect 27663 10013 27675 10047
rect 28810 10044 28816 10056
rect 28771 10016 28816 10044
rect 27617 10007 27675 10013
rect 12897 9979 12955 9985
rect 12897 9976 12909 9979
rect 2746 9948 11560 9976
rect 12406 9948 12909 9976
rect 1394 9868 1400 9920
rect 1452 9908 1458 9920
rect 1949 9911 2007 9917
rect 1949 9908 1961 9911
rect 1452 9880 1961 9908
rect 1452 9868 1458 9880
rect 1949 9877 1961 9880
rect 1995 9877 2007 9911
rect 8938 9908 8944 9920
rect 8899 9880 8944 9908
rect 1949 9871 2007 9877
rect 8938 9868 8944 9880
rect 8996 9868 9002 9920
rect 9030 9868 9036 9920
rect 9088 9908 9094 9920
rect 11149 9911 11207 9917
rect 11149 9908 11161 9911
rect 9088 9880 11161 9908
rect 9088 9868 9094 9880
rect 11149 9877 11161 9880
rect 11195 9908 11207 9911
rect 11238 9908 11244 9920
rect 11195 9880 11244 9908
rect 11195 9877 11207 9880
rect 11149 9871 11207 9877
rect 11238 9868 11244 9880
rect 11296 9868 11302 9920
rect 11532 9908 11560 9948
rect 12897 9945 12909 9948
rect 12943 9945 12955 9979
rect 12897 9939 12955 9945
rect 15194 9936 15200 9988
rect 15252 9976 15258 9988
rect 16022 9976 16028 9988
rect 15252 9948 16028 9976
rect 15252 9936 15258 9948
rect 16022 9936 16028 9948
rect 16080 9936 16086 9988
rect 16209 9979 16267 9985
rect 16209 9945 16221 9979
rect 16255 9945 16267 9979
rect 16390 9976 16396 9988
rect 16351 9948 16396 9976
rect 16209 9939 16267 9945
rect 15010 9908 15016 9920
rect 11532 9880 15016 9908
rect 15010 9868 15016 9880
rect 15068 9868 15074 9920
rect 16224 9908 16252 9939
rect 16390 9936 16396 9948
rect 16448 9936 16454 9988
rect 17494 9985 17500 9988
rect 17488 9939 17500 9985
rect 17552 9976 17558 9988
rect 20800 9979 20858 9985
rect 17552 9948 17588 9976
rect 17494 9936 17500 9939
rect 17552 9936 17558 9948
rect 20800 9945 20812 9979
rect 20846 9976 20858 9979
rect 20898 9976 20904 9988
rect 20846 9948 20904 9976
rect 20846 9945 20858 9948
rect 20800 9939 20858 9945
rect 20898 9936 20904 9948
rect 20956 9936 20962 9988
rect 25860 9979 25918 9985
rect 25860 9945 25872 9979
rect 25906 9976 25918 9979
rect 26142 9976 26148 9988
rect 25906 9948 26148 9976
rect 25906 9945 25918 9948
rect 25860 9939 25918 9945
rect 26142 9936 26148 9948
rect 26200 9936 26206 9988
rect 27632 9976 27660 10007
rect 28810 10004 28816 10016
rect 28868 10004 28874 10056
rect 28997 10047 29055 10053
rect 28997 10013 29009 10047
rect 29043 10013 29055 10047
rect 28997 10007 29055 10013
rect 29012 9976 29040 10007
rect 30466 10004 30472 10056
rect 30524 10044 30530 10056
rect 30837 10047 30895 10053
rect 30837 10044 30849 10047
rect 30524 10016 30849 10044
rect 30524 10004 30530 10016
rect 30837 10013 30849 10016
rect 30883 10013 30895 10047
rect 30837 10007 30895 10013
rect 31021 10047 31079 10053
rect 31021 10013 31033 10047
rect 31067 10044 31079 10047
rect 32030 10044 32036 10056
rect 31067 10016 32036 10044
rect 31067 10013 31079 10016
rect 31021 10007 31079 10013
rect 31036 9976 31064 10007
rect 32030 10004 32036 10016
rect 32088 10004 32094 10056
rect 32232 10053 32260 10084
rect 32217 10047 32275 10053
rect 32217 10013 32229 10047
rect 32263 10013 32275 10047
rect 32217 10007 32275 10013
rect 32582 10004 32588 10056
rect 32640 10044 32646 10056
rect 32677 10047 32735 10053
rect 32677 10044 32689 10047
rect 32640 10016 32689 10044
rect 32640 10004 32646 10016
rect 32677 10013 32689 10016
rect 32723 10013 32735 10047
rect 32784 10044 32812 10084
rect 33778 10044 33784 10056
rect 32784 10016 33784 10044
rect 32677 10007 32735 10013
rect 33778 10004 33784 10016
rect 33836 10004 33842 10056
rect 32922 9979 32980 9985
rect 32922 9976 32934 9979
rect 26344 9948 31064 9976
rect 32048 9948 32934 9976
rect 26344 9920 26372 9948
rect 16758 9908 16764 9920
rect 16224 9880 16764 9908
rect 16758 9868 16764 9880
rect 16816 9868 16822 9920
rect 20714 9868 20720 9920
rect 20772 9908 20778 9920
rect 21726 9908 21732 9920
rect 20772 9880 21732 9908
rect 20772 9868 20778 9880
rect 21726 9868 21732 9880
rect 21784 9908 21790 9920
rect 21913 9911 21971 9917
rect 21913 9908 21925 9911
rect 21784 9880 21925 9908
rect 21784 9868 21790 9880
rect 21913 9877 21925 9880
rect 21959 9877 21971 9911
rect 21913 9871 21971 9877
rect 24949 9911 25007 9917
rect 24949 9877 24961 9911
rect 24995 9908 25007 9911
rect 26326 9908 26332 9920
rect 24995 9880 26332 9908
rect 24995 9877 25007 9880
rect 24949 9871 25007 9877
rect 26326 9868 26332 9880
rect 26384 9868 26390 9920
rect 28902 9908 28908 9920
rect 28863 9880 28908 9908
rect 28902 9868 28908 9880
rect 28960 9868 28966 9920
rect 32048 9917 32076 9948
rect 32922 9945 32934 9948
rect 32968 9945 32980 9979
rect 32922 9939 32980 9945
rect 32033 9911 32091 9917
rect 32033 9877 32045 9911
rect 32079 9877 32091 9911
rect 32033 9871 32091 9877
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 17494 9704 17500 9716
rect 17455 9676 17500 9704
rect 17494 9664 17500 9676
rect 17552 9664 17558 9716
rect 20898 9704 20904 9716
rect 20859 9676 20904 9704
rect 20898 9664 20904 9676
rect 20956 9664 20962 9716
rect 22094 9704 22100 9716
rect 21928 9676 22100 9704
rect 8196 9639 8254 9645
rect 8196 9605 8208 9639
rect 8242 9636 8254 9639
rect 8938 9636 8944 9648
rect 8242 9608 8944 9636
rect 8242 9605 8254 9608
rect 8196 9599 8254 9605
rect 8938 9596 8944 9608
rect 8996 9596 9002 9648
rect 12434 9596 12440 9648
rect 12492 9636 12498 9648
rect 15197 9639 15255 9645
rect 12492 9608 15148 9636
rect 12492 9596 12498 9608
rect 10321 9571 10379 9577
rect 10321 9537 10333 9571
rect 10367 9568 10379 9571
rect 11054 9568 11060 9580
rect 10367 9540 11060 9568
rect 10367 9537 10379 9540
rect 10321 9531 10379 9537
rect 11054 9528 11060 9540
rect 11112 9528 11118 9580
rect 11974 9568 11980 9580
rect 11935 9540 11980 9568
rect 11974 9528 11980 9540
rect 12032 9528 12038 9580
rect 12618 9528 12624 9580
rect 12676 9568 12682 9580
rect 13081 9571 13139 9577
rect 13081 9568 13093 9571
rect 12676 9540 13093 9568
rect 12676 9528 12682 9540
rect 13081 9537 13093 9540
rect 13127 9537 13139 9571
rect 13538 9568 13544 9580
rect 13081 9531 13139 9537
rect 13188 9540 13544 9568
rect 7926 9500 7932 9512
rect 7887 9472 7932 9500
rect 7926 9460 7932 9472
rect 7984 9460 7990 9512
rect 12710 9460 12716 9512
rect 12768 9500 12774 9512
rect 13188 9500 13216 9540
rect 13538 9528 13544 9540
rect 13596 9568 13602 9580
rect 15013 9571 15071 9577
rect 15013 9568 15025 9571
rect 13596 9540 15025 9568
rect 13596 9528 13602 9540
rect 15013 9537 15025 9540
rect 15059 9537 15071 9571
rect 15120 9568 15148 9608
rect 15197 9605 15209 9639
rect 15243 9636 15255 9639
rect 15746 9636 15752 9648
rect 15243 9608 15752 9636
rect 15243 9605 15255 9608
rect 15197 9599 15255 9605
rect 15746 9596 15752 9608
rect 15804 9596 15810 9648
rect 19797 9639 19855 9645
rect 19797 9636 19809 9639
rect 16960 9608 19809 9636
rect 16960 9580 16988 9608
rect 19797 9605 19809 9608
rect 19843 9636 19855 9639
rect 20162 9636 20168 9648
rect 19843 9608 20168 9636
rect 19843 9605 19855 9608
rect 19797 9599 19855 9605
rect 20162 9596 20168 9608
rect 20220 9596 20226 9648
rect 20622 9596 20628 9648
rect 20680 9636 20686 9648
rect 21928 9636 21956 9676
rect 22094 9664 22100 9676
rect 22152 9664 22158 9716
rect 25314 9704 25320 9716
rect 25275 9676 25320 9704
rect 25314 9664 25320 9676
rect 25372 9664 25378 9716
rect 26142 9704 26148 9716
rect 26103 9676 26148 9704
rect 26142 9664 26148 9676
rect 26200 9664 26206 9716
rect 29362 9664 29368 9716
rect 29420 9704 29426 9716
rect 29917 9707 29975 9713
rect 29917 9704 29929 9707
rect 29420 9676 29929 9704
rect 29420 9664 29426 9676
rect 29917 9673 29929 9676
rect 29963 9673 29975 9707
rect 29917 9667 29975 9673
rect 22370 9636 22376 9648
rect 20680 9608 21956 9636
rect 22066 9608 22376 9636
rect 20680 9596 20686 9608
rect 16942 9568 16948 9580
rect 15120 9540 16948 9568
rect 15013 9531 15071 9537
rect 12768 9472 13216 9500
rect 13357 9503 13415 9509
rect 12768 9460 12774 9472
rect 13357 9469 13369 9503
rect 13403 9500 13415 9503
rect 14090 9500 14096 9512
rect 13403 9472 14096 9500
rect 13403 9469 13415 9472
rect 13357 9463 13415 9469
rect 14090 9460 14096 9472
rect 14148 9460 14154 9512
rect 9309 9435 9367 9441
rect 9309 9401 9321 9435
rect 9355 9432 9367 9435
rect 15028 9432 15056 9531
rect 16942 9528 16948 9540
rect 17000 9528 17006 9580
rect 17681 9571 17739 9577
rect 17681 9537 17693 9571
rect 17727 9568 17739 9571
rect 18690 9568 18696 9580
rect 17727 9540 18696 9568
rect 17727 9537 17739 9540
rect 17681 9531 17739 9537
rect 18690 9528 18696 9540
rect 18748 9528 18754 9580
rect 19150 9568 19156 9580
rect 19111 9540 19156 9568
rect 19150 9528 19156 9540
rect 19208 9528 19214 9580
rect 21085 9571 21143 9577
rect 21085 9537 21097 9571
rect 21131 9568 21143 9571
rect 21542 9568 21548 9580
rect 21131 9540 21548 9568
rect 21131 9537 21143 9540
rect 21085 9531 21143 9537
rect 21542 9528 21548 9540
rect 21600 9528 21606 9580
rect 21910 9568 21916 9580
rect 21871 9540 21916 9568
rect 21910 9528 21916 9540
rect 21968 9568 21974 9580
rect 22066 9568 22094 9608
rect 22370 9596 22376 9608
rect 22428 9596 22434 9648
rect 23198 9596 23204 9648
rect 23256 9636 23262 9648
rect 25225 9639 25283 9645
rect 25225 9636 25237 9639
rect 23256 9608 25237 9636
rect 23256 9596 23262 9608
rect 25225 9605 25237 9608
rect 25271 9605 25283 9639
rect 25225 9599 25283 9605
rect 25866 9596 25872 9648
rect 25924 9636 25930 9648
rect 28804 9639 28862 9645
rect 25924 9608 27200 9636
rect 25924 9596 25930 9608
rect 21968 9540 22094 9568
rect 22180 9571 22238 9577
rect 21968 9528 21974 9540
rect 22180 9537 22192 9571
rect 22226 9568 22238 9571
rect 22738 9568 22744 9580
rect 22226 9540 22744 9568
rect 22226 9537 22238 9540
rect 22180 9531 22238 9537
rect 22738 9528 22744 9540
rect 22796 9528 22802 9580
rect 24489 9571 24547 9577
rect 24489 9537 24501 9571
rect 24535 9568 24547 9571
rect 24946 9568 24952 9580
rect 24535 9540 24952 9568
rect 24535 9537 24547 9540
rect 24489 9531 24547 9537
rect 24946 9528 24952 9540
rect 25004 9528 25010 9580
rect 26053 9571 26111 9577
rect 26053 9537 26065 9571
rect 26099 9537 26111 9571
rect 26053 9531 26111 9537
rect 26237 9571 26295 9577
rect 26237 9537 26249 9571
rect 26283 9568 26295 9571
rect 26326 9568 26332 9580
rect 26283 9540 26332 9568
rect 26283 9537 26295 9540
rect 26237 9531 26295 9537
rect 23106 9460 23112 9512
rect 23164 9500 23170 9512
rect 24305 9503 24363 9509
rect 24305 9500 24317 9503
rect 23164 9472 24317 9500
rect 23164 9460 23170 9472
rect 24305 9469 24317 9472
rect 24351 9500 24363 9503
rect 25406 9500 25412 9512
rect 24351 9472 25412 9500
rect 24351 9469 24363 9472
rect 24305 9463 24363 9469
rect 25406 9460 25412 9472
rect 25464 9460 25470 9512
rect 15654 9432 15660 9444
rect 9355 9404 13400 9432
rect 15028 9404 15660 9432
rect 9355 9401 9367 9404
rect 9309 9395 9367 9401
rect 8202 9324 8208 9376
rect 8260 9364 8266 9376
rect 9324 9364 9352 9395
rect 13372 9376 13400 9404
rect 15654 9392 15660 9404
rect 15712 9392 15718 9444
rect 16022 9392 16028 9444
rect 16080 9432 16086 9444
rect 19981 9435 20039 9441
rect 19981 9432 19993 9435
rect 16080 9404 19993 9432
rect 16080 9392 16086 9404
rect 19981 9401 19993 9404
rect 20027 9401 20039 9435
rect 19981 9395 20039 9401
rect 10134 9364 10140 9376
rect 8260 9336 9352 9364
rect 10095 9336 10140 9364
rect 8260 9324 8266 9336
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 11790 9364 11796 9376
rect 11751 9336 11796 9364
rect 11790 9324 11796 9336
rect 11848 9324 11854 9376
rect 12897 9367 12955 9373
rect 12897 9333 12909 9367
rect 12943 9364 12955 9367
rect 12986 9364 12992 9376
rect 12943 9336 12992 9364
rect 12943 9333 12955 9336
rect 12897 9327 12955 9333
rect 12986 9324 12992 9336
rect 13044 9324 13050 9376
rect 13262 9364 13268 9376
rect 13223 9336 13268 9364
rect 13262 9324 13268 9336
rect 13320 9324 13326 9376
rect 13354 9324 13360 9376
rect 13412 9324 13418 9376
rect 18969 9367 19027 9373
rect 18969 9333 18981 9367
rect 19015 9364 19027 9367
rect 19334 9364 19340 9376
rect 19015 9336 19340 9364
rect 19015 9333 19027 9336
rect 18969 9327 19027 9333
rect 19334 9324 19340 9336
rect 19392 9324 19398 9376
rect 19996 9364 20024 9395
rect 22554 9364 22560 9376
rect 19996 9336 22560 9364
rect 22554 9324 22560 9336
rect 22612 9324 22618 9376
rect 22830 9324 22836 9376
rect 22888 9364 22894 9376
rect 23293 9367 23351 9373
rect 23293 9364 23305 9367
rect 22888 9336 23305 9364
rect 22888 9324 22894 9336
rect 23293 9333 23305 9336
rect 23339 9333 23351 9367
rect 23293 9327 23351 9333
rect 24673 9367 24731 9373
rect 24673 9333 24685 9367
rect 24719 9364 24731 9367
rect 25222 9364 25228 9376
rect 24719 9336 25228 9364
rect 24719 9333 24731 9336
rect 24673 9327 24731 9333
rect 25222 9324 25228 9336
rect 25280 9324 25286 9376
rect 26068 9364 26096 9531
rect 26326 9528 26332 9540
rect 26384 9528 26390 9580
rect 26970 9568 26976 9580
rect 26931 9540 26976 9568
rect 26970 9528 26976 9540
rect 27028 9528 27034 9580
rect 27172 9509 27200 9608
rect 28804 9605 28816 9639
rect 28850 9636 28862 9639
rect 28902 9636 28908 9648
rect 28850 9608 28908 9636
rect 28850 9605 28862 9608
rect 28804 9599 28862 9605
rect 28902 9596 28908 9608
rect 28960 9596 28966 9648
rect 30374 9596 30380 9648
rect 30432 9636 30438 9648
rect 30837 9639 30895 9645
rect 30837 9636 30849 9639
rect 30432 9608 30849 9636
rect 30432 9596 30438 9608
rect 30837 9605 30849 9608
rect 30883 9605 30895 9639
rect 30837 9599 30895 9605
rect 32030 9596 32036 9648
rect 32088 9636 32094 9648
rect 32088 9608 32352 9636
rect 32088 9596 32094 9608
rect 27341 9571 27399 9577
rect 27341 9537 27353 9571
rect 27387 9537 27399 9571
rect 27341 9531 27399 9537
rect 31205 9571 31263 9577
rect 31205 9537 31217 9571
rect 31251 9568 31263 9571
rect 31846 9568 31852 9580
rect 31251 9540 31852 9568
rect 31251 9537 31263 9540
rect 31205 9531 31263 9537
rect 27157 9503 27215 9509
rect 27157 9469 27169 9503
rect 27203 9469 27215 9503
rect 27157 9463 27215 9469
rect 26602 9392 26608 9444
rect 26660 9432 26666 9444
rect 27356 9432 27384 9531
rect 31846 9528 31852 9540
rect 31904 9528 31910 9580
rect 32324 9577 32352 9608
rect 32125 9571 32183 9577
rect 32125 9537 32137 9571
rect 32171 9537 32183 9571
rect 32125 9531 32183 9537
rect 32309 9571 32367 9577
rect 32309 9537 32321 9571
rect 32355 9537 32367 9571
rect 32309 9531 32367 9537
rect 27522 9460 27528 9512
rect 27580 9500 27586 9512
rect 28537 9503 28595 9509
rect 28537 9500 28549 9503
rect 27580 9472 28549 9500
rect 27580 9460 27586 9472
rect 28537 9469 28549 9472
rect 28583 9469 28595 9503
rect 28537 9463 28595 9469
rect 29546 9460 29552 9512
rect 29604 9500 29610 9512
rect 30282 9500 30288 9512
rect 29604 9472 30288 9500
rect 29604 9460 29610 9472
rect 30282 9460 30288 9472
rect 30340 9500 30346 9512
rect 31021 9503 31079 9509
rect 31021 9500 31033 9503
rect 30340 9472 31033 9500
rect 30340 9460 30346 9472
rect 31021 9469 31033 9472
rect 31067 9469 31079 9503
rect 31021 9463 31079 9469
rect 31110 9460 31116 9512
rect 31168 9500 31174 9512
rect 31168 9472 31213 9500
rect 31168 9460 31174 9472
rect 32140 9432 32168 9531
rect 26660 9404 27384 9432
rect 31036 9404 32168 9432
rect 26660 9392 26666 9404
rect 27157 9367 27215 9373
rect 27157 9364 27169 9367
rect 26068 9336 27169 9364
rect 27157 9333 27169 9336
rect 27203 9333 27215 9367
rect 27157 9327 27215 9333
rect 27246 9324 27252 9376
rect 27304 9364 27310 9376
rect 31036 9373 31064 9404
rect 31021 9367 31079 9373
rect 27304 9336 27349 9364
rect 27304 9324 27310 9336
rect 31021 9333 31033 9367
rect 31067 9333 31079 9367
rect 32214 9364 32220 9376
rect 32175 9336 32220 9364
rect 31021 9327 31079 9333
rect 32214 9324 32220 9336
rect 32272 9324 32278 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 9122 9120 9128 9172
rect 9180 9160 9186 9172
rect 9309 9163 9367 9169
rect 9309 9160 9321 9163
rect 9180 9132 9321 9160
rect 9180 9120 9186 9132
rect 9309 9129 9321 9132
rect 9355 9129 9367 9163
rect 16022 9160 16028 9172
rect 9309 9123 9367 9129
rect 9416 9132 16028 9160
rect 8938 9052 8944 9104
rect 8996 9092 9002 9104
rect 9416 9092 9444 9132
rect 16022 9120 16028 9132
rect 16080 9120 16086 9172
rect 16206 9160 16212 9172
rect 16167 9132 16212 9160
rect 16206 9120 16212 9132
rect 16264 9120 16270 9172
rect 18690 9160 18696 9172
rect 18651 9132 18696 9160
rect 18690 9120 18696 9132
rect 18748 9120 18754 9172
rect 21542 9160 21548 9172
rect 19260 9132 20208 9160
rect 21503 9132 21548 9160
rect 8996 9064 9444 9092
rect 13081 9095 13139 9101
rect 8996 9052 9002 9064
rect 13081 9061 13093 9095
rect 13127 9092 13139 9095
rect 13906 9092 13912 9104
rect 13127 9064 13912 9092
rect 13127 9061 13139 9064
rect 13081 9055 13139 9061
rect 13906 9052 13912 9064
rect 13964 9052 13970 9104
rect 16577 9095 16635 9101
rect 16577 9061 16589 9095
rect 16623 9092 16635 9095
rect 19260 9092 19288 9132
rect 16623 9064 19288 9092
rect 20180 9092 20208 9132
rect 21542 9120 21548 9132
rect 21600 9120 21606 9172
rect 22094 9120 22100 9172
rect 22152 9160 22158 9172
rect 33134 9160 33140 9172
rect 22152 9132 33140 9160
rect 22152 9120 22158 9132
rect 33134 9120 33140 9132
rect 33192 9120 33198 9172
rect 20180 9064 23060 9092
rect 16623 9061 16635 9064
rect 16577 9055 16635 9061
rect 7926 8984 7932 9036
rect 7984 9024 7990 9036
rect 9582 9024 9588 9036
rect 7984 8996 9588 9024
rect 7984 8984 7990 8996
rect 9582 8984 9588 8996
rect 9640 9024 9646 9036
rect 9640 8996 9812 9024
rect 9640 8984 9646 8996
rect 8938 8956 8944 8968
rect 8899 8928 8944 8956
rect 8938 8916 8944 8928
rect 8996 8916 9002 8968
rect 9122 8956 9128 8968
rect 9083 8928 9128 8956
rect 9122 8916 9128 8928
rect 9180 8916 9186 8968
rect 9784 8965 9812 8996
rect 11514 8984 11520 9036
rect 11572 9024 11578 9036
rect 11701 9027 11759 9033
rect 11701 9024 11713 9027
rect 11572 8996 11713 9024
rect 11572 8984 11578 8996
rect 11701 8993 11713 8996
rect 11747 8993 11759 9027
rect 17313 9027 17371 9033
rect 17313 9024 17325 9027
rect 11701 8987 11759 8993
rect 14660 8996 17325 9024
rect 9769 8959 9827 8965
rect 9769 8925 9781 8959
rect 9815 8956 9827 8959
rect 11532 8956 11560 8984
rect 9815 8928 11560 8956
rect 9815 8925 9827 8928
rect 9769 8919 9827 8925
rect 11790 8916 11796 8968
rect 11848 8956 11854 8968
rect 11957 8959 12015 8965
rect 11957 8956 11969 8959
rect 11848 8928 11969 8956
rect 11848 8916 11854 8928
rect 11957 8925 11969 8928
rect 12003 8925 12015 8959
rect 11957 8919 12015 8925
rect 12342 8916 12348 8968
rect 12400 8956 12406 8968
rect 14660 8965 14688 8996
rect 17313 8993 17325 8996
rect 17359 9024 17371 9027
rect 18322 9024 18328 9036
rect 17359 8996 18328 9024
rect 17359 8993 17371 8996
rect 17313 8987 17371 8993
rect 18322 8984 18328 8996
rect 18380 8984 18386 9036
rect 22830 9024 22836 9036
rect 22296 8996 22836 9024
rect 14645 8959 14703 8965
rect 14645 8956 14657 8959
rect 12400 8928 14657 8956
rect 12400 8916 12406 8928
rect 14645 8925 14657 8928
rect 14691 8925 14703 8959
rect 14826 8956 14832 8968
rect 14787 8928 14832 8956
rect 14645 8919 14703 8925
rect 14826 8916 14832 8928
rect 14884 8916 14890 8968
rect 15013 8959 15071 8965
rect 15013 8925 15025 8959
rect 15059 8956 15071 8959
rect 15657 8959 15715 8965
rect 15657 8956 15669 8959
rect 15059 8928 15669 8956
rect 15059 8925 15071 8928
rect 15013 8919 15071 8925
rect 15657 8925 15669 8928
rect 15703 8925 15715 8959
rect 15657 8919 15715 8925
rect 16117 8959 16175 8965
rect 16117 8925 16129 8959
rect 16163 8925 16175 8959
rect 16117 8919 16175 8925
rect 10036 8891 10094 8897
rect 10036 8857 10048 8891
rect 10082 8888 10094 8891
rect 10134 8888 10140 8900
rect 10082 8860 10140 8888
rect 10082 8857 10094 8860
rect 10036 8851 10094 8857
rect 10134 8848 10140 8860
rect 10192 8848 10198 8900
rect 13262 8848 13268 8900
rect 13320 8888 13326 8900
rect 16132 8888 16160 8919
rect 16942 8916 16948 8968
rect 17000 8956 17006 8968
rect 17037 8959 17095 8965
rect 17037 8956 17049 8959
rect 17000 8928 17049 8956
rect 17000 8916 17006 8928
rect 17037 8925 17049 8928
rect 17083 8925 17095 8959
rect 18506 8956 18512 8968
rect 18467 8928 18512 8956
rect 17037 8919 17095 8925
rect 18506 8916 18512 8928
rect 18564 8916 18570 8968
rect 19242 8956 19248 8968
rect 19203 8928 19248 8956
rect 19242 8916 19248 8928
rect 19300 8916 19306 8968
rect 19334 8916 19340 8968
rect 19392 8956 19398 8968
rect 19501 8959 19559 8965
rect 19501 8956 19513 8959
rect 19392 8928 19513 8956
rect 19392 8916 19398 8928
rect 19501 8925 19513 8928
rect 19547 8925 19559 8959
rect 19501 8919 19559 8925
rect 21177 8959 21235 8965
rect 21177 8925 21189 8959
rect 21223 8925 21235 8959
rect 21358 8956 21364 8968
rect 21319 8928 21364 8956
rect 21177 8919 21235 8925
rect 16666 8888 16672 8900
rect 13320 8860 16672 8888
rect 13320 8848 13326 8860
rect 16666 8848 16672 8860
rect 16724 8848 16730 8900
rect 21192 8888 21220 8919
rect 21358 8916 21364 8928
rect 21416 8916 21422 8968
rect 22051 8959 22109 8965
rect 22051 8925 22063 8959
rect 22097 8956 22109 8959
rect 22296 8956 22324 8996
rect 22830 8984 22836 8996
rect 22888 8984 22894 9036
rect 23032 8968 23060 9064
rect 25406 8984 25412 9036
rect 25464 9024 25470 9036
rect 26878 9024 26884 9036
rect 25464 8996 26884 9024
rect 25464 8984 25470 8996
rect 26878 8984 26884 8996
rect 26936 9024 26942 9036
rect 27617 9027 27675 9033
rect 27617 9024 27629 9027
rect 26936 8996 27629 9024
rect 26936 8984 26942 8996
rect 27617 8993 27629 8996
rect 27663 8993 27675 9027
rect 27617 8987 27675 8993
rect 22097 8928 22324 8956
rect 22373 8959 22431 8965
rect 22097 8925 22109 8928
rect 22051 8919 22109 8925
rect 22373 8925 22385 8959
rect 22419 8956 22431 8959
rect 22419 8928 22683 8956
rect 22419 8925 22431 8928
rect 22373 8919 22431 8925
rect 21450 8888 21456 8900
rect 21192 8860 21456 8888
rect 21450 8848 21456 8860
rect 21508 8848 21514 8900
rect 22186 8888 22192 8900
rect 22147 8860 22192 8888
rect 22186 8848 22192 8860
rect 22244 8848 22250 8900
rect 22278 8848 22284 8900
rect 22336 8888 22342 8900
rect 22336 8860 22381 8888
rect 22336 8848 22342 8860
rect 22655 8832 22683 8928
rect 23014 8916 23020 8968
rect 23072 8956 23078 8968
rect 23072 8928 23117 8956
rect 23072 8916 23078 8928
rect 23198 8916 23204 8968
rect 23256 8956 23262 8968
rect 23293 8959 23351 8965
rect 23293 8956 23305 8959
rect 23256 8928 23305 8956
rect 23256 8916 23262 8928
rect 23293 8925 23305 8928
rect 23339 8925 23351 8959
rect 23293 8919 23351 8925
rect 24397 8959 24455 8965
rect 24397 8925 24409 8959
rect 24443 8956 24455 8959
rect 26234 8956 26240 8968
rect 24443 8928 26240 8956
rect 24443 8925 24455 8928
rect 24397 8919 24455 8925
rect 26234 8916 26240 8928
rect 26292 8916 26298 8968
rect 27801 8959 27859 8965
rect 27801 8925 27813 8959
rect 27847 8956 27859 8959
rect 28994 8956 29000 8968
rect 27847 8928 29000 8956
rect 27847 8925 27859 8928
rect 27801 8919 27859 8925
rect 28994 8916 29000 8928
rect 29052 8916 29058 8968
rect 31021 8959 31079 8965
rect 31021 8925 31033 8959
rect 31067 8956 31079 8959
rect 32582 8956 32588 8968
rect 31067 8928 32588 8956
rect 31067 8925 31079 8928
rect 31021 8919 31079 8925
rect 32582 8916 32588 8928
rect 32640 8916 32646 8968
rect 24664 8891 24722 8897
rect 24664 8857 24676 8891
rect 24710 8888 24722 8891
rect 25130 8888 25136 8900
rect 24710 8860 25136 8888
rect 24710 8857 24722 8860
rect 24664 8851 24722 8857
rect 25130 8848 25136 8860
rect 25188 8848 25194 8900
rect 25314 8848 25320 8900
rect 25372 8888 25378 8900
rect 27246 8888 27252 8900
rect 25372 8860 27252 8888
rect 25372 8848 25378 8860
rect 27246 8848 27252 8860
rect 27304 8848 27310 8900
rect 31288 8891 31346 8897
rect 31288 8857 31300 8891
rect 31334 8888 31346 8891
rect 32214 8888 32220 8900
rect 31334 8860 32220 8888
rect 31334 8857 31346 8860
rect 31288 8851 31346 8857
rect 32214 8848 32220 8860
rect 32272 8848 32278 8900
rect 33045 8891 33103 8897
rect 33045 8857 33057 8891
rect 33091 8888 33103 8891
rect 34606 8888 34612 8900
rect 33091 8860 34612 8888
rect 33091 8857 33103 8860
rect 33045 8851 33103 8857
rect 34606 8848 34612 8860
rect 34664 8848 34670 8900
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 9858 8820 9864 8832
rect 9732 8792 9864 8820
rect 9732 8780 9738 8792
rect 9858 8780 9864 8792
rect 9916 8820 9922 8832
rect 11149 8823 11207 8829
rect 11149 8820 11161 8823
rect 9916 8792 11161 8820
rect 9916 8780 9922 8792
rect 11149 8789 11161 8792
rect 11195 8789 11207 8823
rect 15470 8820 15476 8832
rect 15431 8792 15476 8820
rect 11149 8783 11207 8789
rect 15470 8780 15476 8792
rect 15528 8780 15534 8832
rect 18598 8780 18604 8832
rect 18656 8820 18662 8832
rect 20625 8823 20683 8829
rect 20625 8820 20637 8823
rect 18656 8792 20637 8820
rect 18656 8780 18662 8792
rect 20625 8789 20637 8792
rect 20671 8789 20683 8823
rect 20625 8783 20683 8789
rect 22462 8780 22468 8832
rect 22520 8820 22526 8832
rect 22557 8823 22615 8829
rect 22557 8820 22569 8823
rect 22520 8792 22569 8820
rect 22520 8780 22526 8792
rect 22557 8789 22569 8792
rect 22603 8789 22615 8823
rect 22557 8783 22615 8789
rect 22646 8780 22652 8832
rect 22704 8820 22710 8832
rect 24762 8820 24768 8832
rect 22704 8792 24768 8820
rect 22704 8780 22710 8792
rect 24762 8780 24768 8792
rect 24820 8780 24826 8832
rect 24854 8780 24860 8832
rect 24912 8820 24918 8832
rect 25777 8823 25835 8829
rect 25777 8820 25789 8823
rect 24912 8792 25789 8820
rect 24912 8780 24918 8792
rect 25777 8789 25789 8792
rect 25823 8789 25835 8823
rect 25777 8783 25835 8789
rect 26510 8780 26516 8832
rect 26568 8820 26574 8832
rect 27798 8820 27804 8832
rect 26568 8792 27804 8820
rect 26568 8780 26574 8792
rect 27798 8780 27804 8792
rect 27856 8780 27862 8832
rect 27982 8820 27988 8832
rect 27943 8792 27988 8820
rect 27982 8780 27988 8792
rect 28040 8780 28046 8832
rect 30282 8780 30288 8832
rect 30340 8820 30346 8832
rect 32401 8823 32459 8829
rect 32401 8820 32413 8823
rect 30340 8792 32413 8820
rect 30340 8780 30346 8792
rect 32401 8789 32413 8792
rect 32447 8789 32459 8823
rect 32401 8783 32459 8789
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 8757 8619 8815 8625
rect 8757 8585 8769 8619
rect 8803 8616 8815 8619
rect 9122 8616 9128 8628
rect 8803 8588 9128 8616
rect 8803 8585 8815 8588
rect 8757 8579 8815 8585
rect 9122 8576 9128 8588
rect 9180 8576 9186 8628
rect 11514 8616 11520 8628
rect 10980 8588 11520 8616
rect 4614 8508 4620 8560
rect 4672 8548 4678 8560
rect 10980 8557 11008 8588
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 13906 8616 13912 8628
rect 12406 8588 13912 8616
rect 8481 8551 8539 8557
rect 8481 8548 8493 8551
rect 4672 8520 8493 8548
rect 4672 8508 4678 8520
rect 8481 8517 8493 8520
rect 8527 8517 8539 8551
rect 8481 8511 8539 8517
rect 10965 8551 11023 8557
rect 10965 8517 10977 8551
rect 11011 8517 11023 8551
rect 12406 8548 12434 8588
rect 13906 8576 13912 8588
rect 13964 8576 13970 8628
rect 14090 8576 14096 8628
rect 14148 8616 14154 8628
rect 16206 8616 16212 8628
rect 14148 8588 16212 8616
rect 14148 8576 14154 8588
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 17954 8576 17960 8628
rect 18012 8576 18018 8628
rect 18049 8619 18107 8625
rect 18049 8585 18061 8619
rect 18095 8616 18107 8619
rect 18506 8616 18512 8628
rect 18095 8588 18512 8616
rect 18095 8585 18107 8588
rect 18049 8579 18107 8585
rect 18506 8576 18512 8588
rect 18564 8576 18570 8628
rect 19521 8619 19579 8625
rect 19521 8585 19533 8619
rect 19567 8616 19579 8619
rect 20530 8616 20536 8628
rect 19567 8588 20536 8616
rect 19567 8585 19579 8588
rect 19521 8579 19579 8585
rect 20530 8576 20536 8588
rect 20588 8576 20594 8628
rect 24946 8616 24952 8628
rect 24907 8588 24952 8616
rect 24946 8576 24952 8588
rect 25004 8576 25010 8628
rect 25590 8616 25596 8628
rect 25551 8588 25596 8616
rect 25590 8576 25596 8588
rect 25648 8576 25654 8628
rect 13538 8548 13544 8560
rect 10965 8511 11023 8517
rect 11532 8520 12434 8548
rect 12728 8520 13544 8548
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8449 7711 8483
rect 8202 8480 8208 8492
rect 8163 8452 8208 8480
rect 7653 8443 7711 8449
rect 7668 8344 7696 8443
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 8389 8483 8447 8489
rect 8389 8449 8401 8483
rect 8435 8449 8447 8483
rect 8570 8480 8576 8492
rect 8531 8452 8576 8480
rect 8389 8443 8447 8449
rect 8404 8356 8432 8443
rect 8570 8440 8576 8452
rect 8628 8440 8634 8492
rect 8754 8440 8760 8492
rect 8812 8480 8818 8492
rect 9214 8480 9220 8492
rect 8812 8452 9220 8480
rect 8812 8440 8818 8452
rect 9214 8440 9220 8452
rect 9272 8440 9278 8492
rect 11532 8489 11560 8520
rect 11517 8483 11575 8489
rect 11517 8449 11529 8483
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 11701 8483 11759 8489
rect 11701 8449 11713 8483
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 9858 8372 9864 8424
rect 9916 8412 9922 8424
rect 11716 8412 11744 8443
rect 11790 8440 11796 8492
rect 11848 8480 11854 8492
rect 12728 8489 12756 8520
rect 13538 8508 13544 8520
rect 13596 8508 13602 8560
rect 16114 8548 16120 8560
rect 14660 8520 16120 8548
rect 12986 8489 12992 8492
rect 11931 8483 11989 8489
rect 11848 8452 11893 8480
rect 11848 8440 11854 8452
rect 11931 8449 11943 8483
rect 11977 8480 11989 8483
rect 12713 8483 12771 8489
rect 11977 8452 12204 8480
rect 11977 8449 11989 8452
rect 11931 8443 11989 8449
rect 12066 8412 12072 8424
rect 9916 8384 12072 8412
rect 9916 8372 9922 8384
rect 12066 8372 12072 8384
rect 12124 8372 12130 8424
rect 8386 8344 8392 8356
rect 7668 8316 8248 8344
rect 8299 8316 8392 8344
rect 7466 8276 7472 8288
rect 7427 8248 7472 8276
rect 7466 8236 7472 8248
rect 7524 8236 7530 8288
rect 8220 8276 8248 8316
rect 8386 8304 8392 8316
rect 8444 8344 8450 8356
rect 9876 8344 9904 8372
rect 8444 8316 9904 8344
rect 8444 8304 8450 8316
rect 12176 8288 12204 8452
rect 12713 8449 12725 8483
rect 12759 8449 12771 8483
rect 12980 8480 12992 8489
rect 12947 8452 12992 8480
rect 12713 8443 12771 8449
rect 12980 8443 12992 8452
rect 12986 8440 12992 8443
rect 13044 8440 13050 8492
rect 14660 8489 14688 8520
rect 16114 8508 16120 8520
rect 16172 8508 16178 8560
rect 17972 8548 18000 8576
rect 17512 8520 18000 8548
rect 14645 8483 14703 8489
rect 14645 8449 14657 8483
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 14912 8483 14970 8489
rect 14912 8449 14924 8483
rect 14958 8480 14970 8483
rect 15470 8480 15476 8492
rect 14958 8452 15476 8480
rect 14958 8449 14970 8452
rect 14912 8443 14970 8449
rect 15470 8440 15476 8452
rect 15528 8440 15534 8492
rect 17512 8489 17540 8520
rect 18782 8508 18788 8560
rect 18840 8548 18846 8560
rect 22189 8551 22247 8557
rect 18840 8520 18885 8548
rect 18840 8508 18846 8520
rect 22189 8517 22201 8551
rect 22235 8548 22247 8551
rect 23290 8548 23296 8560
rect 22235 8520 23296 8548
rect 22235 8517 22247 8520
rect 22189 8511 22247 8517
rect 23290 8508 23296 8520
rect 23348 8508 23354 8560
rect 23474 8508 23480 8560
rect 23532 8548 23538 8560
rect 24581 8551 24639 8557
rect 24581 8548 24593 8551
rect 23532 8520 24593 8548
rect 23532 8508 23538 8520
rect 24581 8517 24593 8520
rect 24627 8517 24639 8551
rect 24581 8511 24639 8517
rect 24670 8508 24676 8560
rect 24728 8548 24734 8560
rect 27522 8548 27528 8560
rect 24728 8520 24773 8548
rect 26994 8520 27528 8548
rect 24728 8508 24734 8520
rect 17497 8483 17555 8489
rect 17497 8449 17509 8483
rect 17543 8449 17555 8483
rect 17497 8443 17555 8449
rect 17681 8483 17739 8489
rect 17681 8449 17693 8483
rect 17727 8449 17739 8483
rect 17681 8443 17739 8449
rect 15838 8372 15844 8424
rect 15896 8412 15902 8424
rect 17696 8412 17724 8443
rect 17770 8440 17776 8492
rect 17828 8480 17834 8492
rect 17911 8483 17969 8489
rect 17828 8452 17873 8480
rect 17828 8440 17834 8452
rect 17911 8449 17923 8483
rect 17957 8449 17969 8483
rect 17911 8443 17969 8449
rect 18509 8483 18567 8489
rect 18509 8449 18521 8483
rect 18555 8480 18567 8483
rect 18598 8480 18604 8492
rect 18555 8452 18604 8480
rect 18555 8449 18567 8452
rect 18509 8443 18567 8449
rect 15896 8384 17724 8412
rect 17926 8412 17954 8443
rect 18598 8440 18604 8452
rect 18656 8440 18662 8492
rect 18690 8440 18696 8492
rect 18748 8480 18754 8492
rect 18923 8483 18981 8489
rect 18748 8452 18793 8480
rect 18748 8440 18754 8452
rect 18923 8449 18935 8483
rect 18969 8480 18981 8483
rect 19610 8480 19616 8492
rect 18969 8452 19616 8480
rect 18969 8449 18981 8452
rect 18923 8443 18981 8449
rect 19076 8412 19104 8452
rect 19610 8440 19616 8452
rect 19668 8440 19674 8492
rect 19705 8483 19763 8489
rect 19705 8449 19717 8483
rect 19751 8480 19763 8483
rect 21634 8480 21640 8492
rect 19751 8452 21640 8480
rect 19751 8449 19763 8452
rect 19705 8443 19763 8449
rect 21634 8440 21640 8452
rect 21692 8440 21698 8492
rect 21726 8440 21732 8492
rect 21784 8480 21790 8492
rect 22646 8480 22652 8492
rect 21784 8452 22652 8480
rect 21784 8440 21790 8452
rect 22646 8440 22652 8452
rect 22704 8440 22710 8492
rect 24210 8440 24216 8492
rect 24268 8480 24274 8492
rect 24397 8483 24455 8489
rect 24397 8480 24409 8483
rect 24268 8452 24409 8480
rect 24268 8440 24274 8452
rect 24397 8449 24409 8452
rect 24443 8480 24455 8483
rect 24486 8480 24492 8492
rect 24443 8452 24492 8480
rect 24443 8449 24455 8452
rect 24397 8443 24455 8449
rect 24486 8440 24492 8452
rect 24544 8440 24550 8492
rect 24762 8440 24768 8492
rect 24820 8480 24826 8492
rect 25406 8480 25412 8492
rect 24820 8452 24865 8480
rect 25367 8452 25412 8480
rect 24820 8440 24826 8452
rect 25406 8440 25412 8452
rect 25464 8440 25470 8492
rect 26418 8480 26424 8492
rect 26379 8452 26424 8480
rect 26418 8440 26424 8452
rect 26476 8440 26482 8492
rect 26994 8489 27022 8520
rect 27522 8508 27528 8520
rect 27580 8508 27586 8560
rect 27706 8508 27712 8560
rect 27764 8548 27770 8560
rect 27764 8520 34652 8548
rect 27764 8508 27770 8520
rect 34624 8492 34652 8520
rect 26973 8483 27031 8489
rect 26973 8449 26985 8483
rect 27019 8449 27031 8483
rect 27229 8483 27287 8489
rect 27229 8480 27241 8483
rect 26973 8443 27031 8449
rect 27080 8452 27241 8480
rect 20162 8412 20168 8424
rect 17926 8384 19104 8412
rect 20123 8384 20168 8412
rect 15896 8372 15902 8384
rect 15930 8304 15936 8356
rect 15988 8344 15994 8356
rect 16025 8347 16083 8353
rect 16025 8344 16037 8347
rect 15988 8316 16037 8344
rect 15988 8304 15994 8316
rect 16025 8313 16037 8316
rect 16071 8313 16083 8347
rect 17696 8344 17724 8384
rect 20162 8372 20168 8384
rect 20220 8372 20226 8424
rect 20441 8415 20499 8421
rect 20441 8381 20453 8415
rect 20487 8412 20499 8415
rect 21450 8412 21456 8424
rect 20487 8384 21456 8412
rect 20487 8381 20499 8384
rect 20441 8375 20499 8381
rect 21450 8372 21456 8384
rect 21508 8372 21514 8424
rect 22278 8372 22284 8424
rect 22336 8412 22342 8424
rect 27080 8412 27108 8452
rect 27229 8449 27241 8452
rect 27275 8449 27287 8483
rect 27229 8443 27287 8449
rect 27798 8440 27804 8492
rect 27856 8480 27862 8492
rect 29457 8483 29515 8489
rect 29457 8480 29469 8483
rect 27856 8452 29469 8480
rect 27856 8440 27862 8452
rect 29457 8449 29469 8452
rect 29503 8449 29515 8483
rect 29457 8443 29515 8449
rect 29641 8483 29699 8489
rect 29641 8449 29653 8483
rect 29687 8480 29699 8483
rect 30098 8480 30104 8492
rect 29687 8452 30104 8480
rect 29687 8449 29699 8452
rect 29641 8443 29699 8449
rect 22336 8384 24624 8412
rect 22336 8372 22342 8384
rect 18690 8344 18696 8356
rect 17696 8316 18696 8344
rect 16025 8307 16083 8313
rect 18690 8304 18696 8316
rect 18748 8344 18754 8356
rect 21266 8344 21272 8356
rect 18748 8316 21272 8344
rect 18748 8304 18754 8316
rect 21266 8304 21272 8316
rect 21324 8304 21330 8356
rect 22370 8304 22376 8356
rect 22428 8344 22434 8356
rect 23477 8347 23535 8353
rect 23477 8344 23489 8347
rect 22428 8316 23489 8344
rect 22428 8304 22434 8316
rect 23477 8313 23489 8316
rect 23523 8313 23535 8347
rect 23477 8307 23535 8313
rect 9398 8276 9404 8288
rect 8220 8248 9404 8276
rect 9398 8236 9404 8248
rect 9456 8236 9462 8288
rect 11790 8236 11796 8288
rect 11848 8276 11854 8288
rect 12069 8279 12127 8285
rect 12069 8276 12081 8279
rect 11848 8248 12081 8276
rect 11848 8236 11854 8248
rect 12069 8245 12081 8248
rect 12115 8245 12127 8279
rect 12069 8239 12127 8245
rect 12158 8236 12164 8288
rect 12216 8276 12222 8288
rect 14918 8276 14924 8288
rect 12216 8248 14924 8276
rect 12216 8236 12222 8248
rect 14918 8236 14924 8248
rect 14976 8236 14982 8288
rect 15286 8236 15292 8288
rect 15344 8276 15350 8288
rect 15948 8276 15976 8304
rect 15344 8248 15976 8276
rect 15344 8236 15350 8248
rect 18506 8236 18512 8288
rect 18564 8276 18570 8288
rect 19061 8279 19119 8285
rect 19061 8276 19073 8279
rect 18564 8248 19073 8276
rect 18564 8236 18570 8248
rect 19061 8245 19073 8248
rect 19107 8245 19119 8279
rect 19061 8239 19119 8245
rect 21450 8236 21456 8288
rect 21508 8276 21514 8288
rect 22278 8276 22284 8288
rect 21508 8248 22284 8276
rect 21508 8236 21514 8248
rect 22278 8236 22284 8248
rect 22336 8276 22342 8288
rect 23106 8276 23112 8288
rect 22336 8248 23112 8276
rect 22336 8236 22342 8248
rect 23106 8236 23112 8248
rect 23164 8236 23170 8288
rect 24596 8276 24624 8384
rect 26252 8384 27108 8412
rect 29472 8412 29500 8443
rect 30098 8440 30104 8452
rect 30156 8440 30162 8492
rect 32306 8440 32312 8492
rect 32364 8480 32370 8492
rect 32841 8483 32899 8489
rect 32841 8480 32853 8483
rect 32364 8452 32853 8480
rect 32364 8440 32370 8452
rect 32841 8449 32853 8452
rect 32887 8449 32899 8483
rect 34606 8480 34612 8492
rect 34567 8452 34612 8480
rect 32841 8443 32899 8449
rect 34606 8440 34612 8452
rect 34664 8440 34670 8492
rect 34790 8480 34796 8492
rect 34751 8452 34796 8480
rect 34790 8440 34796 8452
rect 34848 8440 34854 8492
rect 30282 8412 30288 8424
rect 29472 8384 30288 8412
rect 26252 8353 26280 8384
rect 30282 8372 30288 8384
rect 30340 8372 30346 8424
rect 32582 8412 32588 8424
rect 32543 8384 32588 8412
rect 32582 8372 32588 8384
rect 32640 8372 32646 8424
rect 26237 8347 26295 8353
rect 26237 8313 26249 8347
rect 26283 8313 26295 8347
rect 28353 8347 28411 8353
rect 28353 8344 28365 8347
rect 26237 8307 26295 8313
rect 27908 8316 28365 8344
rect 25038 8276 25044 8288
rect 24596 8248 25044 8276
rect 25038 8236 25044 8248
rect 25096 8236 25102 8288
rect 26786 8236 26792 8288
rect 26844 8276 26850 8288
rect 27908 8276 27936 8316
rect 28353 8313 28365 8316
rect 28399 8313 28411 8347
rect 33962 8344 33968 8356
rect 33923 8316 33968 8344
rect 28353 8307 28411 8313
rect 33962 8304 33968 8316
rect 34020 8304 34026 8356
rect 29822 8276 29828 8288
rect 26844 8248 27936 8276
rect 29783 8248 29828 8276
rect 26844 8236 26850 8248
rect 29822 8236 29828 8248
rect 29880 8236 29886 8288
rect 29914 8236 29920 8288
rect 29972 8276 29978 8288
rect 33226 8276 33232 8288
rect 29972 8248 33232 8276
rect 29972 8236 29978 8248
rect 33226 8236 33232 8248
rect 33284 8236 33290 8288
rect 34514 8236 34520 8288
rect 34572 8276 34578 8288
rect 34977 8279 35035 8285
rect 34977 8276 34989 8279
rect 34572 8248 34989 8276
rect 34572 8236 34578 8248
rect 34977 8245 34989 8248
rect 35023 8245 35035 8279
rect 34977 8239 35035 8245
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 8202 8072 8208 8084
rect 8163 8044 8208 8072
rect 8202 8032 8208 8044
rect 8260 8032 8266 8084
rect 11054 8072 11060 8084
rect 11015 8044 11060 8072
rect 11054 8032 11060 8044
rect 11112 8032 11118 8084
rect 11974 8072 11980 8084
rect 11935 8044 11980 8072
rect 11974 8032 11980 8044
rect 12032 8032 12038 8084
rect 14826 8032 14832 8084
rect 14884 8072 14890 8084
rect 15013 8075 15071 8081
rect 15013 8072 15025 8075
rect 14884 8044 15025 8072
rect 14884 8032 14890 8044
rect 15013 8041 15025 8044
rect 15059 8041 15071 8075
rect 15013 8035 15071 8041
rect 15654 8032 15660 8084
rect 15712 8072 15718 8084
rect 18693 8075 18751 8081
rect 15712 8044 16804 8072
rect 15712 8032 15718 8044
rect 12158 8004 12164 8016
rect 10060 7976 12164 8004
rect 8570 7896 8576 7948
rect 8628 7936 8634 7948
rect 10060 7936 10088 7976
rect 12158 7964 12164 7976
rect 12216 7964 12222 8016
rect 12986 7964 12992 8016
rect 13044 8004 13050 8016
rect 15562 8004 15568 8016
rect 13044 7976 15568 8004
rect 13044 7964 13050 7976
rect 15562 7964 15568 7976
rect 15620 7964 15626 8016
rect 16666 8004 16672 8016
rect 16627 7976 16672 8004
rect 16666 7964 16672 7976
rect 16724 7964 16730 8016
rect 16776 8004 16804 8044
rect 18693 8041 18705 8075
rect 18739 8072 18751 8075
rect 19150 8072 19156 8084
rect 18739 8044 19156 8072
rect 18739 8041 18751 8044
rect 18693 8035 18751 8041
rect 19150 8032 19156 8044
rect 19208 8032 19214 8084
rect 21177 8075 21235 8081
rect 19260 8044 20760 8072
rect 19260 8004 19288 8044
rect 16776 7976 19288 8004
rect 20732 8004 20760 8044
rect 21177 8041 21189 8075
rect 21223 8072 21235 8075
rect 21358 8072 21364 8084
rect 21223 8044 21364 8072
rect 21223 8041 21235 8044
rect 21177 8035 21235 8041
rect 21358 8032 21364 8044
rect 21416 8032 21422 8084
rect 21637 8075 21695 8081
rect 21637 8041 21649 8075
rect 21683 8072 21695 8075
rect 22738 8072 22744 8084
rect 21683 8044 22744 8072
rect 21683 8041 21695 8044
rect 21637 8035 21695 8041
rect 22738 8032 22744 8044
rect 22796 8032 22802 8084
rect 25130 8072 25136 8084
rect 25091 8044 25136 8072
rect 25130 8032 25136 8044
rect 25188 8032 25194 8084
rect 25700 8044 28488 8072
rect 23385 8007 23443 8013
rect 23385 8004 23397 8007
rect 20732 7976 23397 8004
rect 23385 7973 23397 7976
rect 23431 8004 23443 8007
rect 25700 8004 25728 8044
rect 28460 8004 28488 8044
rect 28626 8032 28632 8084
rect 28684 8072 28690 8084
rect 28905 8075 28963 8081
rect 28905 8072 28917 8075
rect 28684 8044 28917 8072
rect 28684 8032 28690 8044
rect 28905 8041 28917 8044
rect 28951 8041 28963 8075
rect 28905 8035 28963 8041
rect 29178 8032 29184 8084
rect 29236 8072 29242 8084
rect 31297 8075 31355 8081
rect 31297 8072 31309 8075
rect 29236 8044 31309 8072
rect 29236 8032 29242 8044
rect 31297 8041 31309 8044
rect 31343 8041 31355 8075
rect 33045 8075 33103 8081
rect 33045 8072 33057 8075
rect 31297 8035 31355 8041
rect 32232 8044 33057 8072
rect 29914 8004 29920 8016
rect 23431 7976 25728 8004
rect 26436 7976 27568 8004
rect 28460 7976 29920 8004
rect 23431 7973 23443 7976
rect 23385 7967 23443 7973
rect 8628 7908 10088 7936
rect 8628 7896 8634 7908
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7868 6883 7871
rect 7926 7868 7932 7880
rect 6871 7840 7932 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 7926 7828 7932 7840
rect 7984 7828 7990 7880
rect 9674 7868 9680 7880
rect 9635 7840 9680 7868
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 9858 7868 9864 7880
rect 9819 7840 9864 7868
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 10060 7877 10088 7908
rect 10689 7939 10747 7945
rect 10689 7905 10701 7939
rect 10735 7936 10747 7939
rect 11609 7939 11667 7945
rect 11609 7936 11621 7939
rect 10735 7908 11621 7936
rect 10735 7905 10747 7908
rect 10689 7899 10747 7905
rect 11609 7905 11621 7908
rect 11655 7936 11667 7939
rect 12342 7936 12348 7948
rect 11655 7908 12348 7936
rect 11655 7905 11667 7908
rect 11609 7899 11667 7905
rect 12342 7896 12348 7908
rect 12400 7896 12406 7948
rect 15838 7936 15844 7948
rect 14660 7908 15844 7936
rect 10045 7871 10103 7877
rect 10045 7837 10057 7871
rect 10091 7837 10103 7871
rect 10045 7831 10103 7837
rect 10873 7871 10931 7877
rect 10873 7837 10885 7871
rect 10919 7837 10931 7871
rect 11790 7868 11796 7880
rect 11751 7840 11796 7868
rect 10873 7831 10931 7837
rect 7092 7803 7150 7809
rect 7092 7769 7104 7803
rect 7138 7800 7150 7803
rect 7466 7800 7472 7812
rect 7138 7772 7472 7800
rect 7138 7769 7150 7772
rect 7092 7763 7150 7769
rect 7466 7760 7472 7772
rect 7524 7760 7530 7812
rect 9953 7803 10011 7809
rect 9953 7769 9965 7803
rect 9999 7769 10011 7803
rect 10888 7800 10916 7831
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 14660 7877 14688 7908
rect 15838 7896 15844 7908
rect 15896 7896 15902 7948
rect 16206 7896 16212 7948
rect 16264 7936 16270 7948
rect 16301 7939 16359 7945
rect 16301 7936 16313 7939
rect 16264 7908 16313 7936
rect 16264 7896 16270 7908
rect 16301 7905 16313 7908
rect 16347 7905 16359 7939
rect 16301 7899 16359 7905
rect 16761 7939 16819 7945
rect 16761 7905 16773 7939
rect 16807 7936 16819 7939
rect 17954 7936 17960 7948
rect 16807 7908 17960 7936
rect 16807 7905 16819 7908
rect 16761 7899 16819 7905
rect 17954 7896 17960 7908
rect 18012 7896 18018 7948
rect 18322 7936 18328 7948
rect 18283 7908 18328 7936
rect 18322 7896 18328 7908
rect 18380 7896 18386 7948
rect 18874 7896 18880 7948
rect 18932 7936 18938 7948
rect 19150 7936 19156 7948
rect 18932 7908 19156 7936
rect 18932 7896 18938 7908
rect 19150 7896 19156 7908
rect 19208 7896 19214 7948
rect 19610 7896 19616 7948
rect 19668 7936 19674 7948
rect 19889 7939 19947 7945
rect 19889 7936 19901 7939
rect 19668 7908 19901 7936
rect 19668 7896 19674 7908
rect 19889 7905 19901 7908
rect 19935 7936 19947 7939
rect 22649 7939 22707 7945
rect 22649 7936 22661 7939
rect 19935 7908 21036 7936
rect 19935 7905 19947 7908
rect 19889 7899 19947 7905
rect 14461 7871 14519 7877
rect 14461 7837 14473 7871
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 14645 7871 14703 7877
rect 14645 7837 14657 7871
rect 14691 7837 14703 7871
rect 14645 7831 14703 7837
rect 14829 7871 14887 7877
rect 14829 7837 14841 7871
rect 14875 7870 14887 7871
rect 14918 7870 14924 7880
rect 14875 7842 14924 7870
rect 14875 7837 14887 7842
rect 14829 7831 14887 7837
rect 9953 7763 10011 7769
rect 10244 7772 10916 7800
rect 9490 7692 9496 7744
rect 9548 7732 9554 7744
rect 9968 7732 9996 7763
rect 10244 7741 10272 7772
rect 9548 7704 9996 7732
rect 10229 7735 10287 7741
rect 9548 7692 9554 7704
rect 10229 7701 10241 7735
rect 10275 7701 10287 7735
rect 14476 7732 14504 7831
rect 14918 7828 14924 7842
rect 14976 7868 14982 7880
rect 15470 7868 15476 7880
rect 14976 7840 15069 7868
rect 15431 7840 15476 7868
rect 14976 7828 14982 7840
rect 14550 7760 14556 7812
rect 14608 7800 14614 7812
rect 14737 7803 14795 7809
rect 14737 7800 14749 7803
rect 14608 7772 14749 7800
rect 14608 7760 14614 7772
rect 14737 7769 14749 7772
rect 14783 7769 14795 7803
rect 15028 7800 15056 7840
rect 15470 7828 15476 7840
rect 15528 7828 15534 7880
rect 18506 7868 18512 7880
rect 18467 7840 18512 7868
rect 18506 7828 18512 7840
rect 18564 7828 18570 7880
rect 20625 7871 20683 7877
rect 20625 7837 20637 7871
rect 20671 7868 20683 7871
rect 20714 7868 20720 7880
rect 20671 7840 20720 7868
rect 20671 7837 20683 7840
rect 20625 7831 20683 7837
rect 20714 7828 20720 7840
rect 20772 7828 20778 7880
rect 21008 7877 21036 7908
rect 21836 7908 22661 7936
rect 20993 7871 21051 7877
rect 20993 7837 21005 7871
rect 21039 7868 21051 7871
rect 21726 7868 21732 7880
rect 21039 7840 21732 7868
rect 21039 7837 21051 7840
rect 20993 7831 21051 7837
rect 21726 7828 21732 7840
rect 21784 7828 21790 7880
rect 21836 7877 21864 7908
rect 22649 7905 22661 7908
rect 22695 7905 22707 7939
rect 22649 7899 22707 7905
rect 23290 7896 23296 7948
rect 23348 7936 23354 7948
rect 26234 7936 26240 7948
rect 23348 7908 26240 7936
rect 23348 7896 23354 7908
rect 26234 7896 26240 7908
rect 26292 7896 26298 7948
rect 21821 7871 21879 7877
rect 21821 7837 21833 7871
rect 21867 7837 21879 7871
rect 22278 7868 22284 7880
rect 22239 7840 22284 7868
rect 21821 7831 21879 7837
rect 22278 7828 22284 7840
rect 22336 7828 22342 7880
rect 22462 7868 22468 7880
rect 22423 7840 22468 7868
rect 22462 7828 22468 7840
rect 22520 7828 22526 7880
rect 23198 7868 23204 7880
rect 23159 7840 23204 7868
rect 23198 7828 23204 7840
rect 23256 7868 23262 7880
rect 24397 7871 24455 7877
rect 24397 7868 24409 7871
rect 23256 7840 24409 7868
rect 23256 7828 23262 7840
rect 24397 7837 24409 7840
rect 24443 7837 24455 7871
rect 24397 7831 24455 7837
rect 25222 7828 25228 7880
rect 25280 7868 25286 7880
rect 25317 7871 25375 7877
rect 25317 7868 25329 7871
rect 25280 7840 25329 7868
rect 25280 7828 25286 7840
rect 25317 7837 25329 7840
rect 25363 7837 25375 7871
rect 25317 7831 25375 7837
rect 17681 7803 17739 7809
rect 15028 7772 15424 7800
rect 14737 7763 14795 7769
rect 15286 7732 15292 7744
rect 14476 7704 15292 7732
rect 10229 7695 10287 7701
rect 15286 7692 15292 7704
rect 15344 7692 15350 7744
rect 15396 7732 15424 7772
rect 17681 7769 17693 7803
rect 17727 7800 17739 7803
rect 19426 7800 19432 7812
rect 17727 7772 19432 7800
rect 17727 7769 17739 7772
rect 17681 7763 17739 7769
rect 19426 7760 19432 7772
rect 19484 7800 19490 7812
rect 19705 7803 19763 7809
rect 19705 7800 19717 7803
rect 19484 7772 19717 7800
rect 19484 7760 19490 7772
rect 19705 7769 19717 7772
rect 19751 7769 19763 7803
rect 19705 7763 19763 7769
rect 20809 7803 20867 7809
rect 20809 7769 20821 7803
rect 20855 7769 20867 7803
rect 20809 7763 20867 7769
rect 20901 7803 20959 7809
rect 20901 7769 20913 7803
rect 20947 7800 20959 7803
rect 23290 7800 23296 7812
rect 20947 7772 23296 7800
rect 20947 7769 20959 7772
rect 20901 7763 20959 7769
rect 17773 7735 17831 7741
rect 17773 7732 17785 7735
rect 15396 7704 17785 7732
rect 17773 7701 17785 7704
rect 17819 7701 17831 7735
rect 17773 7695 17831 7701
rect 18046 7692 18052 7744
rect 18104 7732 18110 7744
rect 18506 7732 18512 7744
rect 18104 7704 18512 7732
rect 18104 7692 18110 7704
rect 18506 7692 18512 7704
rect 18564 7692 18570 7744
rect 20824 7732 20852 7763
rect 23290 7760 23296 7772
rect 23348 7760 23354 7812
rect 23474 7760 23480 7812
rect 23532 7800 23538 7812
rect 26436 7800 26464 7976
rect 26786 7936 26792 7948
rect 26528 7908 26792 7936
rect 26528 7877 26556 7908
rect 26786 7896 26792 7908
rect 26844 7896 26850 7948
rect 27540 7936 27568 7976
rect 29914 7964 29920 7976
rect 29972 7964 29978 8016
rect 27540 7908 27660 7936
rect 26513 7871 26571 7877
rect 26513 7837 26525 7871
rect 26559 7837 26571 7871
rect 26878 7868 26884 7880
rect 26839 7840 26884 7868
rect 26513 7831 26571 7837
rect 26878 7828 26884 7840
rect 26936 7828 26942 7880
rect 27522 7868 27528 7880
rect 27483 7840 27528 7868
rect 27522 7828 27528 7840
rect 27580 7828 27586 7880
rect 27632 7868 27660 7908
rect 28350 7868 28356 7880
rect 27632 7840 28356 7868
rect 28350 7828 28356 7840
rect 28408 7828 28414 7880
rect 29638 7828 29644 7880
rect 29696 7868 29702 7880
rect 32232 7877 32260 8044
rect 33045 8041 33057 8044
rect 33091 8041 33103 8075
rect 33045 8035 33103 8041
rect 33137 8075 33195 8081
rect 33137 8041 33149 8075
rect 33183 8072 33195 8075
rect 33226 8072 33232 8084
rect 33183 8044 33232 8072
rect 33183 8041 33195 8044
rect 33137 8035 33195 8041
rect 33226 8032 33232 8044
rect 33284 8032 33290 8084
rect 32306 7964 32312 8016
rect 32364 8004 32370 8016
rect 32364 7976 32409 8004
rect 32364 7964 32370 7976
rect 32582 7964 32588 8016
rect 32640 8004 32646 8016
rect 32640 7976 34744 8004
rect 32640 7964 32646 7976
rect 32674 7896 32680 7948
rect 32732 7936 32738 7948
rect 34716 7945 34744 7976
rect 32861 7939 32919 7945
rect 32861 7936 32873 7939
rect 32732 7908 32873 7936
rect 32732 7896 32738 7908
rect 32861 7905 32873 7908
rect 32907 7905 32919 7939
rect 32861 7899 32919 7905
rect 33045 7939 33103 7945
rect 33045 7905 33057 7939
rect 33091 7905 33103 7939
rect 34701 7939 34759 7945
rect 33045 7899 33103 7905
rect 33244 7908 34652 7936
rect 29917 7871 29975 7877
rect 29917 7868 29929 7871
rect 29696 7840 29929 7868
rect 29696 7828 29702 7840
rect 29917 7837 29929 7840
rect 29963 7837 29975 7871
rect 29917 7831 29975 7837
rect 32217 7871 32275 7877
rect 32217 7837 32229 7871
rect 32263 7837 32275 7871
rect 32217 7831 32275 7837
rect 32401 7871 32459 7877
rect 32401 7837 32413 7871
rect 32447 7837 32459 7871
rect 32401 7831 32459 7837
rect 27798 7809 27804 7812
rect 26697 7803 26755 7809
rect 26697 7800 26709 7803
rect 23532 7772 26709 7800
rect 23532 7760 23538 7772
rect 26697 7769 26709 7772
rect 26743 7769 26755 7803
rect 26697 7763 26755 7769
rect 26789 7803 26847 7809
rect 26789 7769 26801 7803
rect 26835 7800 26847 7803
rect 26835 7772 27752 7800
rect 26835 7769 26847 7772
rect 26789 7763 26847 7769
rect 27724 7744 27752 7772
rect 27792 7763 27804 7809
rect 27856 7800 27862 7812
rect 27856 7772 27892 7800
rect 27798 7760 27804 7763
rect 27856 7760 27862 7772
rect 28074 7760 28080 7812
rect 28132 7800 28138 7812
rect 28902 7800 28908 7812
rect 28132 7772 28908 7800
rect 28132 7760 28138 7772
rect 28902 7760 28908 7772
rect 28960 7760 28966 7812
rect 29454 7760 29460 7812
rect 29512 7800 29518 7812
rect 30162 7803 30220 7809
rect 30162 7800 30174 7803
rect 29512 7772 30174 7800
rect 29512 7760 29518 7772
rect 30162 7769 30174 7772
rect 30208 7769 30220 7803
rect 30162 7763 30220 7769
rect 21266 7732 21272 7744
rect 20824 7704 21272 7732
rect 21266 7692 21272 7704
rect 21324 7692 21330 7744
rect 23566 7692 23572 7744
rect 23624 7732 23630 7744
rect 24581 7735 24639 7741
rect 24581 7732 24593 7735
rect 23624 7704 24593 7732
rect 23624 7692 23630 7704
rect 24581 7701 24593 7704
rect 24627 7732 24639 7735
rect 25314 7732 25320 7744
rect 24627 7704 25320 7732
rect 24627 7701 24639 7704
rect 24581 7695 24639 7701
rect 25314 7692 25320 7704
rect 25372 7692 25378 7744
rect 27065 7735 27123 7741
rect 27065 7701 27077 7735
rect 27111 7732 27123 7735
rect 27246 7732 27252 7744
rect 27111 7704 27252 7732
rect 27111 7701 27123 7704
rect 27065 7695 27123 7701
rect 27246 7692 27252 7704
rect 27304 7692 27310 7744
rect 27706 7692 27712 7744
rect 27764 7692 27770 7744
rect 32416 7732 32444 7831
rect 33060 7800 33088 7899
rect 33244 7877 33272 7908
rect 33229 7871 33287 7877
rect 33229 7837 33241 7871
rect 33275 7837 33287 7871
rect 33962 7868 33968 7880
rect 33229 7831 33287 7837
rect 33336 7840 33968 7868
rect 33336 7800 33364 7840
rect 33962 7828 33968 7840
rect 34020 7828 34026 7880
rect 34149 7871 34207 7877
rect 34149 7837 34161 7871
rect 34195 7868 34207 7871
rect 34514 7868 34520 7880
rect 34195 7840 34520 7868
rect 34195 7837 34207 7840
rect 34149 7831 34207 7837
rect 34514 7828 34520 7840
rect 34572 7828 34578 7880
rect 34624 7868 34652 7908
rect 34701 7905 34713 7939
rect 34747 7905 34759 7939
rect 34701 7899 34759 7905
rect 37182 7868 37188 7880
rect 34624 7840 37188 7868
rect 37182 7828 37188 7840
rect 37240 7828 37246 7880
rect 34946 7803 35004 7809
rect 34946 7800 34958 7803
rect 33060 7772 33364 7800
rect 33980 7772 34958 7800
rect 33134 7732 33140 7744
rect 32416 7704 33140 7732
rect 33134 7692 33140 7704
rect 33192 7692 33198 7744
rect 33980 7741 34008 7772
rect 34946 7769 34958 7772
rect 34992 7769 35004 7803
rect 34946 7763 35004 7769
rect 33965 7735 34023 7741
rect 33965 7701 33977 7735
rect 34011 7701 34023 7735
rect 33965 7695 34023 7701
rect 34606 7692 34612 7744
rect 34664 7732 34670 7744
rect 36081 7735 36139 7741
rect 36081 7732 36093 7735
rect 34664 7704 36093 7732
rect 34664 7692 34670 7704
rect 36081 7701 36093 7704
rect 36127 7701 36139 7735
rect 36081 7695 36139 7701
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 8386 7528 8392 7540
rect 8220 7500 8392 7528
rect 8220 7469 8248 7500
rect 8386 7488 8392 7500
rect 8444 7488 8450 7540
rect 9398 7528 9404 7540
rect 9359 7500 9404 7528
rect 9398 7488 9404 7500
rect 9456 7488 9462 7540
rect 14921 7531 14979 7537
rect 14921 7497 14933 7531
rect 14967 7528 14979 7531
rect 15470 7528 15476 7540
rect 14967 7500 15476 7528
rect 14967 7497 14979 7500
rect 14921 7491 14979 7497
rect 15470 7488 15476 7500
rect 15528 7488 15534 7540
rect 18325 7531 18383 7537
rect 18325 7528 18337 7531
rect 18064 7500 18337 7528
rect 8205 7463 8263 7469
rect 8205 7429 8217 7463
rect 8251 7429 8263 7463
rect 8570 7460 8576 7472
rect 8205 7423 8263 7429
rect 8404 7432 8576 7460
rect 8021 7395 8079 7401
rect 8021 7361 8033 7395
rect 8067 7392 8079 7395
rect 8110 7392 8116 7404
rect 8067 7364 8116 7392
rect 8067 7361 8079 7364
rect 8021 7355 8079 7361
rect 8110 7352 8116 7364
rect 8168 7352 8174 7404
rect 8294 7392 8300 7404
rect 8255 7364 8300 7392
rect 8294 7352 8300 7364
rect 8352 7352 8358 7404
rect 8404 7401 8432 7432
rect 8570 7420 8576 7432
rect 8628 7420 8634 7472
rect 12986 7460 12992 7472
rect 12947 7432 12992 7460
rect 12986 7420 12992 7432
rect 13044 7420 13050 7472
rect 13081 7463 13139 7469
rect 13081 7429 13093 7463
rect 13127 7460 13139 7463
rect 15657 7463 15715 7469
rect 15657 7460 15669 7463
rect 13127 7432 15669 7460
rect 13127 7429 13139 7432
rect 13081 7423 13139 7429
rect 15657 7429 15669 7432
rect 15703 7429 15715 7463
rect 18064 7460 18092 7500
rect 18325 7497 18337 7500
rect 18371 7528 18383 7531
rect 18371 7500 33272 7528
rect 18371 7497 18383 7500
rect 18325 7491 18383 7497
rect 19705 7463 19763 7469
rect 19705 7460 19717 7463
rect 15657 7423 15715 7429
rect 17052 7432 18092 7460
rect 18156 7432 19717 7460
rect 8389 7395 8447 7401
rect 8389 7361 8401 7395
rect 8435 7361 8447 7395
rect 9217 7395 9275 7401
rect 9217 7392 9229 7395
rect 8389 7355 8447 7361
rect 8588 7364 9229 7392
rect 8588 7265 8616 7364
rect 9217 7361 9229 7364
rect 9263 7361 9275 7395
rect 12710 7392 12716 7404
rect 12671 7364 12716 7392
rect 9217 7355 9275 7361
rect 12710 7352 12716 7364
rect 12768 7352 12774 7404
rect 8938 7284 8944 7336
rect 8996 7324 9002 7336
rect 9033 7327 9091 7333
rect 9033 7324 9045 7327
rect 8996 7296 9045 7324
rect 8996 7284 9002 7296
rect 9033 7293 9045 7296
rect 9079 7293 9091 7327
rect 9033 7287 9091 7293
rect 11054 7284 11060 7336
rect 11112 7324 11118 7336
rect 12621 7327 12679 7333
rect 12621 7324 12633 7327
rect 11112 7296 12633 7324
rect 11112 7284 11118 7296
rect 12621 7293 12633 7296
rect 12667 7293 12679 7327
rect 12621 7287 12679 7293
rect 8573 7259 8631 7265
rect 8573 7225 8585 7259
rect 8619 7225 8631 7259
rect 8573 7219 8631 7225
rect 12066 7216 12072 7268
rect 12124 7256 12130 7268
rect 13096 7256 13124 7423
rect 13446 7352 13452 7404
rect 13504 7392 13510 7404
rect 13797 7395 13855 7401
rect 13797 7392 13809 7395
rect 13504 7364 13809 7392
rect 13504 7352 13510 7364
rect 13797 7361 13809 7364
rect 13843 7361 13855 7395
rect 13797 7355 13855 7361
rect 15473 7395 15531 7401
rect 15473 7361 15485 7395
rect 15519 7392 15531 7395
rect 17052 7392 17080 7432
rect 15519 7364 17080 7392
rect 17129 7395 17187 7401
rect 15519 7361 15531 7364
rect 15473 7355 15531 7361
rect 17129 7361 17141 7395
rect 17175 7392 17187 7395
rect 17218 7392 17224 7404
rect 17175 7364 17224 7392
rect 17175 7361 17187 7364
rect 17129 7355 17187 7361
rect 17218 7352 17224 7364
rect 17276 7352 17282 7404
rect 18046 7352 18052 7404
rect 18104 7392 18110 7404
rect 18156 7401 18184 7432
rect 19705 7429 19717 7432
rect 19751 7429 19763 7463
rect 21266 7460 21272 7472
rect 21227 7432 21272 7460
rect 19705 7423 19763 7429
rect 21266 7420 21272 7432
rect 21324 7420 21330 7472
rect 21910 7420 21916 7472
rect 21968 7460 21974 7472
rect 23109 7463 23167 7469
rect 23109 7460 23121 7463
rect 21968 7432 23121 7460
rect 21968 7420 21974 7432
rect 23109 7429 23121 7432
rect 23155 7429 23167 7463
rect 23109 7423 23167 7429
rect 23293 7463 23351 7469
rect 23293 7429 23305 7463
rect 23339 7460 23351 7463
rect 23474 7460 23480 7472
rect 23339 7432 23480 7460
rect 23339 7429 23351 7432
rect 23293 7423 23351 7429
rect 23474 7420 23480 7432
rect 23532 7420 23538 7472
rect 23845 7463 23903 7469
rect 23845 7429 23857 7463
rect 23891 7460 23903 7463
rect 24854 7460 24860 7472
rect 23891 7432 24860 7460
rect 23891 7429 23903 7432
rect 23845 7423 23903 7429
rect 24854 7420 24860 7432
rect 24912 7460 24918 7472
rect 25406 7460 25412 7472
rect 24912 7432 25412 7460
rect 24912 7420 24918 7432
rect 25406 7420 25412 7432
rect 25464 7420 25470 7472
rect 26418 7420 26424 7472
rect 26476 7460 26482 7472
rect 27341 7463 27399 7469
rect 27341 7460 27353 7463
rect 26476 7432 27353 7460
rect 26476 7420 26482 7432
rect 27341 7429 27353 7432
rect 27387 7429 27399 7463
rect 27341 7423 27399 7429
rect 28350 7420 28356 7472
rect 28408 7460 28414 7472
rect 28629 7463 28687 7469
rect 28629 7460 28641 7463
rect 28408 7432 28641 7460
rect 28408 7420 28414 7432
rect 28629 7429 28641 7432
rect 28675 7429 28687 7463
rect 28629 7423 28687 7429
rect 28721 7463 28779 7469
rect 28721 7429 28733 7463
rect 28767 7460 28779 7463
rect 30006 7460 30012 7472
rect 28767 7432 30012 7460
rect 28767 7429 28779 7432
rect 28721 7423 28779 7429
rect 30006 7420 30012 7432
rect 30064 7420 30070 7472
rect 33134 7420 33140 7472
rect 33192 7420 33198 7472
rect 33244 7460 33272 7500
rect 34790 7488 34796 7540
rect 34848 7528 34854 7540
rect 35161 7531 35219 7537
rect 35161 7528 35173 7531
rect 34848 7500 35173 7528
rect 34848 7488 34854 7500
rect 35161 7497 35173 7500
rect 35207 7497 35219 7531
rect 35161 7491 35219 7497
rect 34330 7460 34336 7472
rect 33244 7432 34336 7460
rect 34330 7420 34336 7432
rect 34388 7460 34394 7472
rect 34885 7463 34943 7469
rect 34388 7432 34836 7460
rect 34388 7420 34394 7432
rect 18141 7395 18199 7401
rect 18141 7392 18153 7395
rect 18104 7364 18153 7392
rect 18104 7352 18110 7364
rect 18141 7361 18153 7364
rect 18187 7361 18199 7395
rect 18141 7355 18199 7361
rect 18969 7395 19027 7401
rect 18969 7361 18981 7395
rect 19015 7361 19027 7395
rect 20530 7392 20536 7404
rect 20491 7364 20536 7392
rect 18969 7355 19027 7361
rect 13538 7324 13544 7336
rect 13499 7296 13544 7324
rect 13538 7284 13544 7296
rect 13596 7284 13602 7336
rect 17954 7284 17960 7336
rect 18012 7324 18018 7336
rect 18984 7324 19012 7355
rect 20530 7352 20536 7364
rect 20588 7352 20594 7404
rect 21085 7395 21143 7401
rect 21085 7361 21097 7395
rect 21131 7392 21143 7395
rect 21928 7392 21956 7420
rect 21131 7364 21956 7392
rect 22373 7395 22431 7401
rect 21131 7361 21143 7364
rect 21085 7355 21143 7361
rect 22373 7361 22385 7395
rect 22419 7392 22431 7395
rect 22462 7392 22468 7404
rect 22419 7364 22468 7392
rect 22419 7361 22431 7364
rect 22373 7355 22431 7361
rect 18012 7296 19012 7324
rect 19889 7327 19947 7333
rect 18012 7284 18018 7296
rect 19889 7293 19901 7327
rect 19935 7324 19947 7327
rect 21100 7324 21128 7355
rect 22462 7352 22468 7364
rect 22520 7352 22526 7404
rect 23014 7352 23020 7404
rect 23072 7392 23078 7404
rect 23753 7395 23811 7401
rect 23753 7392 23765 7395
rect 23072 7364 23765 7392
rect 23072 7352 23078 7364
rect 23753 7361 23765 7364
rect 23799 7361 23811 7395
rect 23934 7392 23940 7404
rect 23895 7364 23940 7392
rect 23753 7355 23811 7361
rect 23934 7352 23940 7364
rect 23992 7352 23998 7404
rect 26326 7392 26332 7404
rect 26287 7364 26332 7392
rect 26326 7352 26332 7364
rect 26384 7352 26390 7404
rect 26878 7352 26884 7404
rect 26936 7392 26942 7404
rect 27157 7395 27215 7401
rect 26936 7364 27108 7392
rect 26936 7352 26942 7364
rect 19935 7296 21128 7324
rect 19935 7293 19947 7296
rect 19889 7287 19947 7293
rect 22002 7284 22008 7336
rect 22060 7324 22066 7336
rect 22189 7327 22247 7333
rect 22189 7324 22201 7327
rect 22060 7296 22201 7324
rect 22060 7284 22066 7296
rect 22189 7293 22201 7296
rect 22235 7293 22247 7327
rect 22189 7287 22247 7293
rect 24857 7327 24915 7333
rect 24857 7293 24869 7327
rect 24903 7324 24915 7327
rect 24946 7324 24952 7336
rect 24903 7296 24952 7324
rect 24903 7293 24915 7296
rect 24857 7287 24915 7293
rect 24946 7284 24952 7296
rect 25004 7284 25010 7336
rect 25130 7324 25136 7336
rect 25091 7296 25136 7324
rect 25130 7284 25136 7296
rect 25188 7284 25194 7336
rect 26970 7324 26976 7336
rect 26931 7296 26976 7324
rect 26970 7284 26976 7296
rect 27028 7284 27034 7336
rect 27080 7324 27108 7364
rect 27157 7361 27169 7395
rect 27203 7392 27215 7395
rect 27246 7392 27252 7404
rect 27203 7364 27252 7392
rect 27203 7361 27215 7364
rect 27157 7355 27215 7361
rect 27246 7352 27252 7364
rect 27304 7352 27310 7404
rect 27982 7392 27988 7404
rect 27943 7364 27988 7392
rect 27982 7352 27988 7364
rect 28040 7352 28046 7404
rect 28445 7395 28503 7401
rect 28445 7361 28457 7395
rect 28491 7392 28503 7395
rect 28534 7392 28540 7404
rect 28491 7364 28540 7392
rect 28491 7361 28503 7364
rect 28445 7355 28503 7361
rect 28534 7352 28540 7364
rect 28592 7352 28598 7404
rect 28813 7395 28871 7401
rect 28813 7361 28825 7395
rect 28859 7361 28871 7395
rect 28813 7355 28871 7361
rect 29641 7395 29699 7401
rect 29641 7361 29653 7395
rect 29687 7392 29699 7395
rect 29822 7392 29828 7404
rect 29687 7364 29828 7392
rect 29687 7361 29699 7364
rect 29641 7355 29699 7361
rect 28828 7324 28856 7355
rect 29822 7352 29828 7364
rect 29880 7352 29886 7404
rect 30374 7401 30380 7404
rect 30368 7355 30380 7401
rect 30432 7392 30438 7404
rect 32585 7395 32643 7401
rect 30432 7364 30468 7392
rect 30374 7352 30380 7355
rect 30432 7352 30438 7364
rect 32585 7361 32597 7395
rect 32631 7361 32643 7395
rect 32585 7355 32643 7361
rect 32769 7395 32827 7401
rect 32769 7361 32781 7395
rect 32815 7392 32827 7395
rect 33152 7392 33180 7420
rect 34606 7392 34612 7404
rect 32815 7364 33180 7392
rect 34567 7364 34612 7392
rect 32815 7361 32827 7364
rect 32769 7355 32827 7361
rect 27080 7296 28856 7324
rect 30101 7327 30159 7333
rect 30101 7293 30113 7327
rect 30147 7293 30159 7327
rect 32600 7324 32628 7355
rect 34606 7352 34612 7364
rect 34664 7352 34670 7404
rect 34808 7401 34836 7432
rect 34885 7429 34897 7463
rect 34931 7460 34943 7463
rect 37918 7460 37924 7472
rect 34931 7432 37924 7460
rect 34931 7429 34943 7432
rect 34885 7423 34943 7429
rect 37918 7420 37924 7432
rect 37976 7420 37982 7472
rect 34793 7395 34851 7401
rect 34793 7361 34805 7395
rect 34839 7361 34851 7395
rect 34793 7355 34851 7361
rect 34977 7395 35035 7401
rect 34977 7361 34989 7395
rect 35023 7361 35035 7395
rect 34977 7355 35035 7361
rect 33134 7324 33140 7336
rect 32600 7296 33140 7324
rect 30101 7287 30159 7293
rect 12124 7228 13124 7256
rect 19153 7259 19211 7265
rect 12124 7216 12130 7228
rect 19153 7225 19165 7259
rect 19199 7256 19211 7259
rect 19199 7228 19334 7256
rect 19199 7225 19211 7228
rect 19153 7219 19211 7225
rect 12437 7191 12495 7197
rect 12437 7157 12449 7191
rect 12483 7188 12495 7191
rect 13354 7188 13360 7200
rect 12483 7160 13360 7188
rect 12483 7157 12495 7160
rect 12437 7151 12495 7157
rect 13354 7148 13360 7160
rect 13412 7148 13418 7200
rect 16666 7148 16672 7200
rect 16724 7188 16730 7200
rect 17221 7191 17279 7197
rect 17221 7188 17233 7191
rect 16724 7160 17233 7188
rect 16724 7148 16730 7160
rect 17221 7157 17233 7160
rect 17267 7157 17279 7191
rect 19306 7188 19334 7228
rect 19426 7216 19432 7268
rect 19484 7256 19490 7268
rect 19484 7228 29592 7256
rect 19484 7216 19490 7228
rect 19518 7188 19524 7200
rect 19306 7160 19524 7188
rect 17221 7151 17279 7157
rect 19518 7148 19524 7160
rect 19576 7148 19582 7200
rect 20346 7188 20352 7200
rect 20307 7160 20352 7188
rect 20346 7148 20352 7160
rect 20404 7148 20410 7200
rect 22557 7191 22615 7197
rect 22557 7157 22569 7191
rect 22603 7188 22615 7191
rect 23014 7188 23020 7200
rect 22603 7160 23020 7188
rect 22603 7157 22615 7160
rect 22557 7151 22615 7157
rect 23014 7148 23020 7160
rect 23072 7148 23078 7200
rect 25314 7148 25320 7200
rect 25372 7188 25378 7200
rect 26145 7191 26203 7197
rect 26145 7188 26157 7191
rect 25372 7160 26157 7188
rect 25372 7148 25378 7160
rect 26145 7157 26157 7160
rect 26191 7157 26203 7191
rect 27798 7188 27804 7200
rect 27759 7160 27804 7188
rect 26145 7151 26203 7157
rect 27798 7148 27804 7160
rect 27856 7148 27862 7200
rect 28350 7148 28356 7200
rect 28408 7188 28414 7200
rect 28718 7188 28724 7200
rect 28408 7160 28724 7188
rect 28408 7148 28414 7160
rect 28718 7148 28724 7160
rect 28776 7148 28782 7200
rect 28994 7188 29000 7200
rect 28955 7160 29000 7188
rect 28994 7148 29000 7160
rect 29052 7148 29058 7200
rect 29454 7188 29460 7200
rect 29415 7160 29460 7188
rect 29454 7148 29460 7160
rect 29512 7148 29518 7200
rect 29564 7188 29592 7228
rect 29638 7216 29644 7268
rect 29696 7256 29702 7268
rect 30116 7256 30144 7287
rect 33134 7284 33140 7296
rect 33192 7284 33198 7336
rect 34992 7256 35020 7355
rect 35434 7256 35440 7268
rect 29696 7228 30144 7256
rect 31036 7228 35440 7256
rect 29696 7216 29702 7228
rect 31036 7188 31064 7228
rect 35434 7216 35440 7228
rect 35492 7216 35498 7268
rect 31478 7188 31484 7200
rect 29564 7160 31064 7188
rect 31439 7160 31484 7188
rect 31478 7148 31484 7160
rect 31536 7148 31542 7200
rect 32674 7188 32680 7200
rect 32635 7160 32680 7188
rect 32674 7148 32680 7160
rect 32732 7148 32738 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 18046 6984 18052 6996
rect 18007 6956 18052 6984
rect 18046 6944 18052 6956
rect 18104 6944 18110 6996
rect 19426 6944 19432 6996
rect 19484 6984 19490 6996
rect 19705 6987 19763 6993
rect 19705 6984 19717 6987
rect 19484 6956 19717 6984
rect 19484 6944 19490 6956
rect 19705 6953 19717 6956
rect 19751 6953 19763 6987
rect 19705 6947 19763 6953
rect 20272 6956 21312 6984
rect 9582 6808 9588 6860
rect 9640 6848 9646 6860
rect 9861 6851 9919 6857
rect 9861 6848 9873 6851
rect 9640 6820 9873 6848
rect 9640 6808 9646 6820
rect 9861 6817 9873 6820
rect 9907 6817 9919 6851
rect 12986 6848 12992 6860
rect 9861 6811 9919 6817
rect 11716 6820 12992 6848
rect 8938 6740 8944 6792
rect 8996 6780 9002 6792
rect 9217 6783 9275 6789
rect 9217 6780 9229 6783
rect 8996 6752 9229 6780
rect 8996 6740 9002 6752
rect 9217 6749 9229 6752
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6780 9459 6783
rect 9447 6752 10272 6780
rect 9447 6749 9459 6752
rect 9401 6743 9459 6749
rect 8386 6672 8392 6724
rect 8444 6712 8450 6724
rect 9306 6712 9312 6724
rect 8444 6684 9312 6712
rect 8444 6672 8450 6684
rect 9306 6672 9312 6684
rect 9364 6712 9370 6724
rect 9416 6712 9444 6743
rect 9364 6684 9444 6712
rect 9364 6672 9370 6684
rect 9950 6672 9956 6724
rect 10008 6712 10014 6724
rect 10106 6715 10164 6721
rect 10106 6712 10118 6715
rect 10008 6684 10118 6712
rect 10008 6672 10014 6684
rect 10106 6681 10118 6684
rect 10152 6681 10164 6715
rect 10244 6712 10272 6752
rect 10594 6740 10600 6792
rect 10652 6780 10658 6792
rect 11716 6789 11744 6820
rect 12986 6808 12992 6820
rect 13044 6808 13050 6860
rect 13446 6848 13452 6860
rect 13407 6820 13452 6848
rect 13446 6808 13452 6820
rect 13504 6808 13510 6860
rect 16114 6848 16120 6860
rect 13556 6820 15700 6848
rect 16075 6820 16120 6848
rect 11701 6783 11759 6789
rect 11701 6780 11713 6783
rect 10652 6752 11713 6780
rect 10652 6740 10658 6752
rect 11701 6749 11713 6752
rect 11747 6749 11759 6783
rect 11701 6743 11759 6749
rect 11885 6783 11943 6789
rect 11885 6749 11897 6783
rect 11931 6780 11943 6783
rect 11974 6780 11980 6792
rect 11931 6752 11980 6780
rect 11931 6749 11943 6752
rect 11885 6743 11943 6749
rect 11974 6740 11980 6752
rect 12032 6740 12038 6792
rect 12069 6783 12127 6789
rect 12069 6749 12081 6783
rect 12115 6780 12127 6783
rect 12713 6783 12771 6789
rect 12713 6780 12725 6783
rect 12115 6752 12725 6780
rect 12115 6749 12127 6752
rect 12069 6743 12127 6749
rect 12713 6749 12725 6752
rect 12759 6749 12771 6783
rect 13354 6780 13360 6792
rect 13315 6752 13360 6780
rect 12713 6743 12771 6749
rect 13354 6740 13360 6752
rect 13412 6740 13418 6792
rect 13556 6789 13584 6820
rect 13541 6783 13599 6789
rect 13541 6749 13553 6783
rect 13587 6749 13599 6783
rect 15470 6780 15476 6792
rect 15431 6752 15476 6780
rect 13541 6743 13599 6749
rect 11146 6712 11152 6724
rect 10244 6684 11152 6712
rect 10106 6675 10164 6681
rect 11146 6672 11152 6684
rect 11204 6672 11210 6724
rect 11256 6684 12664 6712
rect 10410 6604 10416 6656
rect 10468 6644 10474 6656
rect 11256 6653 11284 6684
rect 11241 6647 11299 6653
rect 11241 6644 11253 6647
rect 10468 6616 11253 6644
rect 10468 6604 10474 6616
rect 11241 6613 11253 6616
rect 11287 6613 11299 6647
rect 12526 6644 12532 6656
rect 12487 6616 12532 6644
rect 11241 6607 11299 6613
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 12636 6644 12664 6684
rect 12894 6672 12900 6724
rect 12952 6712 12958 6724
rect 13556 6712 13584 6743
rect 15470 6740 15476 6752
rect 15528 6740 15534 6792
rect 15672 6789 15700 6820
rect 16114 6808 16120 6820
rect 16172 6808 16178 6860
rect 18138 6808 18144 6860
rect 18196 6848 18202 6860
rect 20272 6848 20300 6956
rect 21284 6916 21312 6956
rect 21358 6944 21364 6996
rect 21416 6984 21422 6996
rect 22002 6984 22008 6996
rect 21416 6956 22008 6984
rect 21416 6944 21422 6956
rect 22002 6944 22008 6956
rect 22060 6984 22066 6996
rect 25130 6984 25136 6996
rect 22060 6956 25136 6984
rect 22060 6944 22066 6956
rect 25130 6944 25136 6956
rect 25188 6984 25194 6996
rect 26418 6984 26424 6996
rect 25188 6956 26424 6984
rect 25188 6944 25194 6956
rect 26418 6944 26424 6956
rect 26476 6944 26482 6996
rect 26970 6944 26976 6996
rect 27028 6984 27034 6996
rect 27522 6984 27528 6996
rect 27028 6956 27528 6984
rect 27028 6944 27034 6956
rect 27522 6944 27528 6956
rect 27580 6984 27586 6996
rect 27709 6987 27767 6993
rect 27709 6984 27721 6987
rect 27580 6956 27721 6984
rect 27580 6944 27586 6956
rect 27709 6953 27721 6956
rect 27755 6953 27767 6987
rect 27709 6947 27767 6953
rect 28994 6944 29000 6996
rect 29052 6984 29058 6996
rect 31478 6984 31484 6996
rect 29052 6956 31484 6984
rect 29052 6944 29058 6956
rect 31478 6944 31484 6956
rect 31536 6944 31542 6996
rect 33962 6944 33968 6996
rect 34020 6984 34026 6996
rect 34701 6987 34759 6993
rect 34701 6984 34713 6987
rect 34020 6956 34713 6984
rect 34020 6944 34026 6956
rect 34701 6953 34713 6956
rect 34747 6953 34759 6987
rect 34701 6947 34759 6953
rect 21637 6919 21695 6925
rect 21637 6916 21649 6919
rect 21284 6888 21649 6916
rect 21637 6885 21649 6888
rect 21683 6885 21695 6919
rect 21637 6879 21695 6885
rect 24670 6876 24676 6928
rect 24728 6916 24734 6928
rect 28074 6916 28080 6928
rect 24728 6888 28080 6916
rect 24728 6876 24734 6888
rect 28074 6876 28080 6888
rect 28132 6876 28138 6928
rect 22370 6848 22376 6860
rect 18196 6820 20300 6848
rect 22066 6820 22376 6848
rect 18196 6808 18202 6820
rect 22066 6792 22094 6820
rect 22370 6808 22376 6820
rect 22428 6808 22434 6860
rect 24118 6808 24124 6860
rect 24176 6848 24182 6860
rect 32306 6848 32312 6860
rect 24176 6820 25912 6848
rect 24176 6808 24182 6820
rect 15657 6783 15715 6789
rect 15657 6749 15669 6783
rect 15703 6749 15715 6783
rect 15657 6743 15715 6749
rect 17954 6740 17960 6792
rect 18012 6780 18018 6792
rect 18049 6783 18107 6789
rect 18049 6780 18061 6783
rect 18012 6752 18061 6780
rect 18012 6740 18018 6752
rect 18049 6749 18061 6752
rect 18095 6749 18107 6783
rect 18230 6780 18236 6792
rect 18191 6752 18236 6780
rect 18049 6743 18107 6749
rect 18230 6740 18236 6752
rect 18288 6740 18294 6792
rect 19518 6780 19524 6792
rect 19479 6752 19524 6780
rect 19518 6740 19524 6752
rect 19576 6740 19582 6792
rect 20257 6783 20315 6789
rect 20257 6749 20269 6783
rect 20303 6780 20315 6783
rect 22066 6780 22100 6792
rect 20303 6752 22100 6780
rect 20303 6749 20315 6752
rect 20257 6743 20315 6749
rect 22094 6740 22100 6752
rect 22152 6740 22158 6792
rect 22278 6740 22284 6792
rect 22336 6780 22342 6792
rect 24581 6783 24639 6789
rect 24581 6780 24593 6783
rect 22336 6752 24593 6780
rect 22336 6740 22342 6752
rect 24581 6749 24593 6752
rect 24627 6749 24639 6783
rect 24581 6743 24639 6749
rect 24670 6740 24676 6792
rect 24728 6780 24734 6792
rect 25884 6789 25912 6820
rect 26436 6820 32312 6848
rect 25225 6783 25283 6789
rect 25225 6780 25237 6783
rect 24728 6752 25237 6780
rect 24728 6740 24734 6752
rect 25225 6749 25237 6752
rect 25271 6749 25283 6783
rect 25225 6743 25283 6749
rect 25869 6783 25927 6789
rect 25869 6749 25881 6783
rect 25915 6749 25927 6783
rect 25869 6743 25927 6749
rect 26234 6740 26240 6792
rect 26292 6780 26298 6792
rect 26436 6789 26464 6820
rect 32306 6808 32312 6820
rect 32364 6808 32370 6860
rect 34885 6851 34943 6857
rect 34885 6817 34897 6851
rect 34931 6848 34943 6851
rect 35802 6848 35808 6860
rect 34931 6820 35808 6848
rect 34931 6817 34943 6820
rect 34885 6811 34943 6817
rect 35802 6808 35808 6820
rect 35860 6808 35866 6860
rect 26421 6783 26479 6789
rect 26421 6780 26433 6783
rect 26292 6752 26433 6780
rect 26292 6740 26298 6752
rect 26421 6749 26433 6752
rect 26467 6749 26479 6783
rect 28813 6783 28871 6789
rect 28813 6780 28825 6783
rect 26421 6743 26479 6749
rect 26528 6752 28825 6780
rect 12952 6684 13584 6712
rect 15565 6715 15623 6721
rect 12952 6672 12958 6684
rect 15565 6681 15577 6715
rect 15611 6712 15623 6715
rect 16362 6715 16420 6721
rect 16362 6712 16374 6715
rect 15611 6684 16374 6712
rect 15611 6681 15623 6684
rect 15565 6675 15623 6681
rect 16362 6681 16374 6684
rect 16408 6681 16420 6715
rect 16362 6675 16420 6681
rect 17512 6684 19840 6712
rect 14274 6644 14280 6656
rect 12636 6616 14280 6644
rect 14274 6604 14280 6616
rect 14332 6604 14338 6656
rect 16850 6604 16856 6656
rect 16908 6644 16914 6656
rect 17512 6653 17540 6684
rect 17497 6647 17555 6653
rect 17497 6644 17509 6647
rect 16908 6616 17509 6644
rect 16908 6604 16914 6616
rect 17497 6613 17509 6616
rect 17543 6613 17555 6647
rect 19812 6644 19840 6684
rect 20346 6672 20352 6724
rect 20404 6712 20410 6724
rect 20502 6715 20560 6721
rect 20502 6712 20514 6715
rect 20404 6684 20514 6712
rect 20404 6672 20410 6684
rect 20502 6681 20514 6684
rect 20548 6681 20560 6715
rect 20502 6675 20560 6681
rect 22640 6715 22698 6721
rect 22640 6681 22652 6715
rect 22686 6712 22698 6715
rect 22830 6712 22836 6724
rect 22686 6684 22836 6712
rect 22686 6681 22698 6684
rect 22640 6675 22698 6681
rect 22830 6672 22836 6684
rect 22888 6672 22894 6724
rect 23290 6672 23296 6724
rect 23348 6712 23354 6724
rect 23348 6684 24440 6712
rect 23348 6672 23354 6684
rect 20622 6644 20628 6656
rect 19812 6616 20628 6644
rect 17497 6607 17555 6613
rect 20622 6604 20628 6616
rect 20680 6604 20686 6656
rect 21818 6604 21824 6656
rect 21876 6644 21882 6656
rect 22186 6644 22192 6656
rect 21876 6616 22192 6644
rect 21876 6604 21882 6616
rect 22186 6604 22192 6616
rect 22244 6644 22250 6656
rect 24412 6653 24440 6684
rect 24486 6672 24492 6724
rect 24544 6712 24550 6724
rect 24544 6684 25728 6712
rect 24544 6672 24550 6684
rect 23753 6647 23811 6653
rect 23753 6644 23765 6647
rect 22244 6616 23765 6644
rect 22244 6604 22250 6616
rect 23753 6613 23765 6616
rect 23799 6613 23811 6647
rect 23753 6607 23811 6613
rect 24397 6647 24455 6653
rect 24397 6613 24409 6647
rect 24443 6613 24455 6647
rect 25038 6644 25044 6656
rect 24999 6616 25044 6644
rect 24397 6607 24455 6613
rect 25038 6604 25044 6616
rect 25096 6604 25102 6656
rect 25700 6653 25728 6684
rect 26050 6672 26056 6724
rect 26108 6712 26114 6724
rect 26528 6712 26556 6752
rect 28813 6749 28825 6752
rect 28859 6749 28871 6783
rect 28813 6743 28871 6749
rect 29178 6740 29184 6792
rect 29236 6780 29242 6792
rect 29549 6783 29607 6789
rect 29549 6780 29561 6783
rect 29236 6752 29561 6780
rect 29236 6740 29242 6752
rect 29549 6749 29561 6752
rect 29595 6749 29607 6783
rect 29914 6780 29920 6792
rect 29875 6752 29920 6780
rect 29549 6743 29607 6749
rect 29914 6740 29920 6752
rect 29972 6740 29978 6792
rect 30282 6740 30288 6792
rect 30340 6780 30346 6792
rect 30561 6783 30619 6789
rect 30561 6780 30573 6783
rect 30340 6752 30573 6780
rect 30340 6740 30346 6752
rect 30561 6749 30573 6752
rect 30607 6749 30619 6783
rect 30742 6780 30748 6792
rect 30703 6752 30748 6780
rect 30561 6743 30619 6749
rect 30742 6740 30748 6752
rect 30800 6740 30806 6792
rect 31754 6740 31760 6792
rect 31812 6780 31818 6792
rect 31812 6752 31857 6780
rect 31812 6740 31818 6752
rect 32122 6740 32128 6792
rect 32180 6780 32186 6792
rect 32674 6789 32680 6792
rect 32401 6783 32459 6789
rect 32401 6780 32413 6783
rect 32180 6752 32413 6780
rect 32180 6740 32186 6752
rect 32401 6749 32413 6752
rect 32447 6749 32459 6783
rect 32668 6780 32680 6789
rect 32635 6752 32680 6780
rect 32401 6743 32459 6749
rect 32668 6743 32680 6752
rect 32674 6740 32680 6743
rect 32732 6740 32738 6792
rect 34606 6740 34612 6792
rect 34664 6780 34670 6792
rect 34977 6783 35035 6789
rect 34977 6780 34989 6783
rect 34664 6752 34989 6780
rect 34664 6740 34670 6752
rect 34977 6749 34989 6752
rect 35023 6749 35035 6783
rect 34977 6743 35035 6749
rect 26108 6684 26556 6712
rect 26108 6672 26114 6684
rect 27614 6672 27620 6724
rect 27672 6712 27678 6724
rect 27672 6684 28672 6712
rect 27672 6672 27678 6684
rect 28644 6653 28672 6684
rect 28718 6672 28724 6724
rect 28776 6712 28782 6724
rect 29270 6712 29276 6724
rect 28776 6684 29276 6712
rect 28776 6672 28782 6684
rect 29270 6672 29276 6684
rect 29328 6712 29334 6724
rect 29733 6715 29791 6721
rect 29733 6712 29745 6715
rect 29328 6684 29745 6712
rect 29328 6672 29334 6684
rect 29733 6681 29745 6684
rect 29779 6681 29791 6715
rect 29733 6675 29791 6681
rect 29825 6715 29883 6721
rect 29825 6681 29837 6715
rect 29871 6712 29883 6715
rect 34701 6715 34759 6721
rect 34701 6712 34713 6715
rect 29871 6684 31616 6712
rect 29871 6681 29883 6684
rect 29825 6675 29883 6681
rect 25685 6647 25743 6653
rect 25685 6613 25697 6647
rect 25731 6613 25743 6647
rect 25685 6607 25743 6613
rect 28629 6647 28687 6653
rect 28629 6613 28641 6647
rect 28675 6613 28687 6647
rect 30098 6644 30104 6656
rect 30059 6616 30104 6644
rect 28629 6607 28687 6613
rect 30098 6604 30104 6616
rect 30156 6604 30162 6656
rect 30466 6604 30472 6656
rect 30524 6644 30530 6656
rect 31588 6653 31616 6684
rect 33796 6684 34713 6712
rect 30929 6647 30987 6653
rect 30929 6644 30941 6647
rect 30524 6616 30941 6644
rect 30524 6604 30530 6616
rect 30929 6613 30941 6616
rect 30975 6613 30987 6647
rect 30929 6607 30987 6613
rect 31573 6647 31631 6653
rect 31573 6613 31585 6647
rect 31619 6613 31631 6647
rect 31573 6607 31631 6613
rect 33318 6604 33324 6656
rect 33376 6644 33382 6656
rect 33796 6653 33824 6684
rect 34701 6681 34713 6684
rect 34747 6681 34759 6715
rect 34701 6675 34759 6681
rect 33781 6647 33839 6653
rect 33781 6644 33793 6647
rect 33376 6616 33793 6644
rect 33376 6604 33382 6616
rect 33781 6613 33793 6616
rect 33827 6613 33839 6647
rect 33781 6607 33839 6613
rect 34790 6604 34796 6656
rect 34848 6644 34854 6656
rect 35161 6647 35219 6653
rect 35161 6644 35173 6647
rect 34848 6616 35173 6644
rect 34848 6604 34854 6616
rect 35161 6613 35173 6616
rect 35207 6613 35219 6647
rect 35161 6607 35219 6613
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 8386 6440 8392 6452
rect 7944 6412 8392 6440
rect 7742 6304 7748 6316
rect 7703 6276 7748 6304
rect 7742 6264 7748 6276
rect 7800 6264 7806 6316
rect 7944 6313 7972 6412
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 9122 6400 9128 6452
rect 9180 6440 9186 6452
rect 9769 6443 9827 6449
rect 9769 6440 9781 6443
rect 9180 6412 9781 6440
rect 9180 6400 9186 6412
rect 9769 6409 9781 6412
rect 9815 6440 9827 6443
rect 9815 6412 13124 6440
rect 9815 6409 9827 6412
rect 9769 6403 9827 6409
rect 8478 6372 8484 6384
rect 8391 6344 8484 6372
rect 8404 6313 8432 6344
rect 8478 6332 8484 6344
rect 8536 6372 8542 6384
rect 9582 6372 9588 6384
rect 8536 6344 9588 6372
rect 8536 6332 8542 6344
rect 9582 6332 9588 6344
rect 9640 6332 9646 6384
rect 10686 6372 10692 6384
rect 10647 6344 10692 6372
rect 10686 6332 10692 6344
rect 10744 6332 10750 6384
rect 11968 6375 12026 6381
rect 11968 6341 11980 6375
rect 12014 6372 12026 6375
rect 12526 6372 12532 6384
rect 12014 6344 12532 6372
rect 12014 6341 12026 6344
rect 11968 6335 12026 6341
rect 12526 6332 12532 6344
rect 12584 6332 12590 6384
rect 13096 6372 13124 6412
rect 13170 6400 13176 6452
rect 13228 6440 13234 6452
rect 13541 6443 13599 6449
rect 13541 6440 13553 6443
rect 13228 6412 13553 6440
rect 13228 6400 13234 6412
rect 13541 6409 13553 6412
rect 13587 6409 13599 6443
rect 13541 6403 13599 6409
rect 14185 6443 14243 6449
rect 14185 6409 14197 6443
rect 14231 6440 14243 6443
rect 14550 6440 14556 6452
rect 14231 6412 14556 6440
rect 14231 6409 14243 6412
rect 14185 6403 14243 6409
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 15102 6440 15108 6452
rect 15063 6412 15108 6440
rect 15102 6400 15108 6412
rect 15160 6400 15166 6452
rect 17497 6443 17555 6449
rect 15212 6412 16896 6440
rect 13814 6372 13820 6384
rect 13096 6344 13820 6372
rect 13814 6332 13820 6344
rect 13872 6332 13878 6384
rect 15212 6372 15240 6412
rect 13924 6344 15240 6372
rect 7929 6307 7987 6313
rect 7929 6273 7941 6307
rect 7975 6273 7987 6307
rect 7929 6267 7987 6273
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6273 8447 6307
rect 8645 6307 8703 6313
rect 8645 6304 8657 6307
rect 8389 6267 8447 6273
rect 8496 6276 8657 6304
rect 7837 6239 7895 6245
rect 7837 6205 7849 6239
rect 7883 6236 7895 6239
rect 8496 6236 8524 6276
rect 8645 6273 8657 6276
rect 8691 6273 8703 6307
rect 10410 6304 10416 6316
rect 10371 6276 10416 6304
rect 8645 6267 8703 6273
rect 10410 6264 10416 6276
rect 10468 6264 10474 6316
rect 10597 6307 10655 6313
rect 10597 6273 10609 6307
rect 10643 6273 10655 6307
rect 10597 6267 10655 6273
rect 10781 6307 10839 6313
rect 10781 6273 10793 6307
rect 10827 6304 10839 6307
rect 11790 6304 11796 6316
rect 10827 6276 11796 6304
rect 10827 6273 10839 6276
rect 10781 6267 10839 6273
rect 7883 6208 8524 6236
rect 10612 6236 10640 6267
rect 11790 6264 11796 6276
rect 11848 6264 11854 6316
rect 12894 6264 12900 6316
rect 12952 6304 12958 6316
rect 13725 6307 13783 6313
rect 13725 6304 13737 6307
rect 12952 6276 13737 6304
rect 12952 6264 12958 6276
rect 13725 6273 13737 6276
rect 13771 6273 13783 6307
rect 13725 6267 13783 6273
rect 11606 6236 11612 6248
rect 10612 6208 11612 6236
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 11606 6196 11612 6208
rect 11664 6196 11670 6248
rect 11701 6239 11759 6245
rect 11701 6205 11713 6239
rect 11747 6205 11759 6239
rect 11701 6199 11759 6205
rect 10778 6060 10784 6112
rect 10836 6100 10842 6112
rect 10965 6103 11023 6109
rect 10965 6100 10977 6103
rect 10836 6072 10977 6100
rect 10836 6060 10842 6072
rect 10965 6069 10977 6072
rect 11011 6069 11023 6103
rect 11716 6100 11744 6199
rect 12802 6196 12808 6248
rect 12860 6236 12866 6248
rect 13924 6236 13952 6344
rect 15470 6332 15476 6384
rect 15528 6372 15534 6384
rect 16739 6375 16797 6381
rect 16739 6372 16751 6375
rect 15528 6344 16751 6372
rect 15528 6332 15534 6344
rect 16739 6341 16751 6344
rect 16785 6341 16797 6375
rect 16868 6372 16896 6412
rect 17497 6409 17509 6443
rect 17543 6440 17555 6443
rect 17586 6440 17592 6452
rect 17543 6412 17592 6440
rect 17543 6409 17555 6412
rect 17497 6403 17555 6409
rect 17586 6400 17592 6412
rect 17644 6400 17650 6452
rect 18598 6440 18604 6452
rect 17696 6412 18604 6440
rect 17696 6372 17724 6412
rect 18598 6400 18604 6412
rect 18656 6400 18662 6452
rect 18690 6400 18696 6452
rect 18748 6440 18754 6452
rect 20162 6440 20168 6452
rect 18748 6412 20168 6440
rect 18748 6400 18754 6412
rect 20162 6400 20168 6412
rect 20220 6400 20226 6452
rect 20349 6443 20407 6449
rect 20349 6409 20361 6443
rect 20395 6440 20407 6443
rect 20530 6440 20536 6452
rect 20395 6412 20536 6440
rect 20395 6409 20407 6412
rect 20349 6403 20407 6409
rect 20530 6400 20536 6412
rect 20588 6400 20594 6452
rect 20622 6400 20628 6452
rect 20680 6440 20686 6452
rect 22373 6443 22431 6449
rect 20680 6412 22324 6440
rect 20680 6400 20686 6412
rect 16868 6344 17724 6372
rect 16739 6335 16797 6341
rect 18138 6332 18144 6384
rect 18196 6372 18202 6384
rect 18785 6375 18843 6381
rect 18785 6372 18797 6375
rect 18196 6344 18797 6372
rect 18196 6332 18202 6344
rect 18785 6341 18797 6344
rect 18831 6341 18843 6375
rect 21358 6372 21364 6384
rect 18785 6335 18843 6341
rect 20088 6344 21364 6372
rect 14090 6264 14096 6316
rect 14148 6304 14154 6316
rect 14369 6307 14427 6313
rect 14369 6304 14381 6307
rect 14148 6276 14381 6304
rect 14148 6264 14154 6276
rect 14369 6273 14381 6276
rect 14415 6273 14427 6307
rect 14369 6267 14427 6273
rect 15010 6264 15016 6316
rect 15068 6304 15074 6316
rect 15289 6307 15347 6313
rect 15289 6304 15301 6307
rect 15068 6276 15301 6304
rect 15068 6264 15074 6276
rect 15289 6273 15301 6276
rect 15335 6273 15347 6307
rect 17037 6307 17095 6313
rect 15289 6267 15347 6273
rect 15396 6276 16988 6304
rect 12860 6208 13952 6236
rect 12860 6196 12866 6208
rect 14734 6196 14740 6248
rect 14792 6236 14798 6248
rect 15396 6236 15424 6276
rect 16666 6236 16672 6248
rect 14792 6208 15424 6236
rect 16627 6208 16672 6236
rect 14792 6196 14798 6208
rect 16666 6196 16672 6208
rect 16724 6196 16730 6248
rect 16850 6236 16856 6248
rect 16811 6208 16856 6236
rect 16850 6196 16856 6208
rect 16908 6196 16914 6248
rect 16960 6236 16988 6276
rect 17037 6273 17049 6307
rect 17083 6304 17095 6307
rect 17126 6304 17132 6316
rect 17083 6276 17132 6304
rect 17083 6273 17095 6276
rect 17037 6267 17095 6273
rect 17126 6264 17132 6276
rect 17184 6264 17190 6316
rect 17402 6264 17408 6316
rect 17460 6304 17466 6316
rect 17681 6307 17739 6313
rect 17681 6304 17693 6307
rect 17460 6276 17693 6304
rect 17460 6264 17466 6276
rect 17681 6273 17693 6276
rect 17727 6273 17739 6307
rect 17681 6267 17739 6273
rect 18230 6264 18236 6316
rect 18288 6304 18294 6316
rect 18509 6307 18567 6313
rect 18509 6304 18521 6307
rect 18288 6276 18521 6304
rect 18288 6264 18294 6276
rect 18509 6273 18521 6276
rect 18555 6273 18567 6307
rect 18690 6304 18696 6316
rect 18651 6276 18696 6304
rect 18509 6267 18567 6273
rect 18690 6264 18696 6276
rect 18748 6264 18754 6316
rect 20088 6313 20116 6344
rect 21358 6332 21364 6344
rect 21416 6332 21422 6384
rect 22296 6372 22324 6412
rect 22373 6409 22385 6443
rect 22419 6440 22431 6443
rect 22462 6440 22468 6452
rect 22419 6412 22468 6440
rect 22419 6409 22431 6412
rect 22373 6403 22431 6409
rect 22462 6400 22468 6412
rect 22520 6400 22526 6452
rect 22830 6440 22836 6452
rect 22791 6412 22836 6440
rect 22830 6400 22836 6412
rect 22888 6400 22894 6452
rect 24489 6443 24547 6449
rect 24489 6409 24501 6443
rect 24535 6440 24547 6443
rect 26234 6440 26240 6452
rect 24535 6412 26240 6440
rect 24535 6409 24547 6412
rect 24489 6403 24547 6409
rect 26234 6400 26240 6412
rect 26292 6400 26298 6452
rect 26421 6443 26479 6449
rect 26421 6409 26433 6443
rect 26467 6440 26479 6443
rect 27062 6440 27068 6452
rect 26467 6412 27068 6440
rect 26467 6409 26479 6412
rect 26421 6403 26479 6409
rect 27062 6400 27068 6412
rect 27120 6400 27126 6452
rect 28074 6440 28080 6452
rect 28035 6412 28080 6440
rect 28074 6400 28080 6412
rect 28132 6400 28138 6452
rect 29733 6443 29791 6449
rect 29733 6409 29745 6443
rect 29779 6409 29791 6443
rect 29733 6403 29791 6409
rect 30285 6443 30343 6449
rect 30285 6409 30297 6443
rect 30331 6440 30343 6443
rect 30374 6440 30380 6452
rect 30331 6412 30380 6440
rect 30331 6409 30343 6412
rect 30285 6403 30343 6409
rect 22922 6372 22928 6384
rect 21468 6344 22232 6372
rect 22296 6344 22928 6372
rect 18877 6307 18935 6313
rect 18877 6273 18889 6307
rect 18923 6273 18935 6307
rect 18877 6267 18935 6273
rect 20073 6307 20131 6313
rect 20073 6273 20085 6307
rect 20119 6273 20131 6307
rect 20073 6267 20131 6273
rect 20165 6307 20223 6313
rect 20165 6273 20177 6307
rect 20211 6304 20223 6307
rect 21082 6304 21088 6316
rect 20211 6276 20300 6304
rect 21043 6276 21088 6304
rect 20211 6273 20223 6276
rect 20165 6267 20223 6273
rect 17310 6236 17316 6248
rect 16960 6208 17316 6236
rect 17310 6196 17316 6208
rect 17368 6196 17374 6248
rect 18598 6196 18604 6248
rect 18656 6236 18662 6248
rect 18892 6236 18920 6267
rect 18656 6208 19012 6236
rect 18656 6196 18662 6208
rect 14182 6128 14188 6180
rect 14240 6168 14246 6180
rect 16684 6168 16712 6196
rect 16942 6168 16948 6180
rect 14240 6140 16712 6168
rect 16903 6140 16948 6168
rect 14240 6128 14246 6140
rect 16942 6128 16948 6140
rect 17000 6168 17006 6180
rect 18874 6168 18880 6180
rect 17000 6140 18880 6168
rect 17000 6128 17006 6140
rect 18874 6128 18880 6140
rect 18932 6128 18938 6180
rect 12434 6100 12440 6112
rect 11716 6072 12440 6100
rect 10965 6063 11023 6069
rect 12434 6060 12440 6072
rect 12492 6060 12498 6112
rect 12710 6060 12716 6112
rect 12768 6100 12774 6112
rect 13081 6103 13139 6109
rect 13081 6100 13093 6103
rect 12768 6072 13093 6100
rect 12768 6060 12774 6072
rect 13081 6069 13093 6072
rect 13127 6100 13139 6103
rect 13906 6100 13912 6112
rect 13127 6072 13912 6100
rect 13127 6069 13139 6072
rect 13081 6063 13139 6069
rect 13906 6060 13912 6072
rect 13964 6060 13970 6112
rect 14642 6060 14648 6112
rect 14700 6100 14706 6112
rect 18690 6100 18696 6112
rect 14700 6072 18696 6100
rect 14700 6060 14706 6072
rect 18690 6060 18696 6072
rect 18748 6060 18754 6112
rect 18984 6100 19012 6208
rect 19061 6171 19119 6177
rect 19061 6137 19073 6171
rect 19107 6168 19119 6171
rect 20272 6168 20300 6276
rect 21082 6264 21088 6276
rect 21140 6264 21146 6316
rect 21468 6304 21496 6344
rect 21818 6304 21824 6316
rect 21192 6276 21496 6304
rect 21779 6276 21824 6304
rect 19107 6140 20300 6168
rect 19107 6137 19119 6140
rect 19061 6131 19119 6137
rect 21192 6109 21220 6276
rect 21818 6264 21824 6276
rect 21876 6264 21882 6316
rect 22204 6313 22232 6344
rect 22922 6332 22928 6344
rect 22980 6332 22986 6384
rect 24397 6375 24455 6381
rect 24397 6341 24409 6375
rect 24443 6372 24455 6375
rect 24854 6372 24860 6384
rect 24443 6344 24860 6372
rect 24443 6341 24455 6344
rect 24397 6335 24455 6341
rect 24854 6332 24860 6344
rect 24912 6332 24918 6384
rect 26970 6372 26976 6384
rect 25056 6344 26976 6372
rect 25056 6316 25084 6344
rect 26970 6332 26976 6344
rect 27028 6332 27034 6384
rect 29748 6372 29776 6403
rect 30374 6400 30380 6412
rect 30432 6400 30438 6452
rect 30929 6443 30987 6449
rect 30929 6409 30941 6443
rect 30975 6440 30987 6443
rect 31018 6440 31024 6452
rect 30975 6412 31024 6440
rect 30975 6409 30987 6412
rect 30929 6403 30987 6409
rect 31018 6400 31024 6412
rect 31076 6400 31082 6452
rect 32232 6412 32536 6440
rect 30742 6372 30748 6384
rect 27448 6344 29592 6372
rect 29748 6344 30748 6372
rect 27448 6316 27476 6344
rect 22005 6307 22063 6313
rect 22005 6273 22017 6307
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 22097 6307 22155 6313
rect 22097 6273 22109 6307
rect 22143 6273 22155 6307
rect 22097 6267 22155 6273
rect 22189 6307 22247 6313
rect 22189 6273 22201 6307
rect 22235 6273 22247 6307
rect 23014 6304 23020 6316
rect 22975 6276 23020 6304
rect 22189 6267 22247 6273
rect 21177 6103 21235 6109
rect 21177 6100 21189 6103
rect 18984 6072 21189 6100
rect 21177 6069 21189 6072
rect 21223 6069 21235 6103
rect 21177 6063 21235 6069
rect 21726 6060 21732 6112
rect 21784 6100 21790 6112
rect 22020 6100 22048 6267
rect 22112 6236 22140 6267
rect 23014 6264 23020 6276
rect 23072 6264 23078 6316
rect 23750 6304 23756 6316
rect 23711 6276 23756 6304
rect 23750 6264 23756 6276
rect 23808 6264 23814 6316
rect 25038 6304 25044 6316
rect 24951 6276 25044 6304
rect 25038 6264 25044 6276
rect 25096 6264 25102 6316
rect 25314 6313 25320 6316
rect 25308 6304 25320 6313
rect 25275 6276 25320 6304
rect 25308 6267 25320 6276
rect 25314 6264 25320 6267
rect 25372 6264 25378 6316
rect 27062 6304 27068 6316
rect 27023 6276 27068 6304
rect 27062 6264 27068 6276
rect 27120 6264 27126 6316
rect 27249 6307 27307 6313
rect 27249 6273 27261 6307
rect 27295 6273 27307 6307
rect 27249 6267 27307 6273
rect 27341 6307 27399 6313
rect 27341 6273 27353 6307
rect 27387 6273 27399 6307
rect 27341 6267 27399 6273
rect 22462 6236 22468 6248
rect 22112 6208 22468 6236
rect 22462 6196 22468 6208
rect 22520 6196 22526 6248
rect 22738 6196 22744 6248
rect 22796 6236 22802 6248
rect 24670 6236 24676 6248
rect 22796 6208 24676 6236
rect 22796 6196 22802 6208
rect 24670 6196 24676 6208
rect 24728 6196 24734 6248
rect 27264 6168 27292 6267
rect 27356 6236 27384 6267
rect 27430 6264 27436 6316
rect 27488 6304 27494 6316
rect 27488 6276 27533 6304
rect 27488 6264 27494 6276
rect 27614 6264 27620 6316
rect 27672 6304 27678 6316
rect 28261 6307 28319 6313
rect 28261 6304 28273 6307
rect 27672 6276 28273 6304
rect 27672 6264 27678 6276
rect 28261 6273 28273 6276
rect 28307 6273 28319 6307
rect 28261 6267 28319 6273
rect 28994 6264 29000 6316
rect 29052 6304 29058 6316
rect 29181 6307 29239 6313
rect 29181 6304 29193 6307
rect 29052 6276 29193 6304
rect 29052 6264 29058 6276
rect 29181 6273 29193 6276
rect 29227 6273 29239 6307
rect 29181 6267 29239 6273
rect 29270 6264 29276 6316
rect 29328 6313 29334 6316
rect 29328 6307 29377 6313
rect 29328 6273 29331 6307
rect 29365 6273 29377 6307
rect 29454 6304 29460 6316
rect 29415 6276 29460 6304
rect 29328 6267 29377 6273
rect 29328 6264 29334 6267
rect 29454 6264 29460 6276
rect 29512 6264 29518 6316
rect 29564 6313 29592 6344
rect 30742 6332 30748 6344
rect 30800 6332 30806 6384
rect 31202 6332 31208 6384
rect 31260 6372 31266 6384
rect 32232 6381 32260 6412
rect 32217 6375 32275 6381
rect 32217 6372 32229 6375
rect 31260 6344 32229 6372
rect 31260 6332 31266 6344
rect 32217 6341 32229 6344
rect 32263 6341 32275 6375
rect 32508 6372 32536 6412
rect 32766 6400 32772 6452
rect 32824 6440 32830 6452
rect 33873 6443 33931 6449
rect 33873 6440 33885 6443
rect 32824 6412 33885 6440
rect 32824 6400 32830 6412
rect 33873 6409 33885 6412
rect 33919 6409 33931 6443
rect 33873 6403 33931 6409
rect 33045 6375 33103 6381
rect 33045 6372 33057 6375
rect 32508 6344 33057 6372
rect 32217 6335 32275 6341
rect 33045 6341 33057 6344
rect 33091 6341 33103 6375
rect 33045 6335 33103 6341
rect 29549 6307 29607 6313
rect 29549 6273 29561 6307
rect 29595 6304 29607 6307
rect 29914 6304 29920 6316
rect 29595 6276 29920 6304
rect 29595 6273 29607 6276
rect 29549 6267 29607 6273
rect 29914 6264 29920 6276
rect 29972 6264 29978 6316
rect 30466 6304 30472 6316
rect 30427 6276 30472 6304
rect 30466 6264 30472 6276
rect 30524 6264 30530 6316
rect 31110 6304 31116 6316
rect 31071 6276 31116 6304
rect 31110 6264 31116 6276
rect 31168 6264 31174 6316
rect 32585 6307 32643 6313
rect 32585 6273 32597 6307
rect 32631 6304 32643 6307
rect 32950 6304 32956 6316
rect 32631 6276 32956 6304
rect 32631 6273 32643 6276
rect 32585 6267 32643 6273
rect 32950 6264 32956 6276
rect 33008 6264 33014 6316
rect 33318 6264 33324 6316
rect 33376 6264 33382 6316
rect 33413 6307 33471 6313
rect 33413 6273 33425 6307
rect 33459 6273 33471 6307
rect 34054 6304 34060 6316
rect 34015 6276 34060 6304
rect 33413 6267 33471 6273
rect 27356 6208 28994 6236
rect 23492 6140 23980 6168
rect 23492 6100 23520 6140
rect 21784 6072 23520 6100
rect 23569 6103 23627 6109
rect 21784 6060 21790 6072
rect 23569 6069 23581 6103
rect 23615 6100 23627 6103
rect 23842 6100 23848 6112
rect 23615 6072 23848 6100
rect 23615 6069 23627 6072
rect 23569 6063 23627 6069
rect 23842 6060 23848 6072
rect 23900 6060 23906 6112
rect 23952 6100 23980 6140
rect 25976 6140 27292 6168
rect 28966 6168 28994 6208
rect 31938 6196 31944 6248
rect 31996 6236 32002 6248
rect 32287 6239 32345 6245
rect 32287 6236 32299 6239
rect 31996 6208 32299 6236
rect 31996 6196 32002 6208
rect 32287 6205 32299 6208
rect 32333 6205 32345 6239
rect 32287 6199 32345 6205
rect 32398 6196 32404 6248
rect 32456 6236 32462 6248
rect 33229 6239 33287 6245
rect 32456 6208 32501 6236
rect 32456 6196 32462 6208
rect 33229 6205 33241 6239
rect 33275 6236 33287 6239
rect 33336 6236 33364 6264
rect 33275 6208 33364 6236
rect 33428 6236 33456 6267
rect 34054 6264 34060 6276
rect 34112 6264 34118 6316
rect 35618 6236 35624 6248
rect 33428 6208 35624 6236
rect 33275 6205 33287 6208
rect 33229 6199 33287 6205
rect 35618 6196 35624 6208
rect 35676 6196 35682 6248
rect 31662 6168 31668 6180
rect 28966 6140 31668 6168
rect 25976 6100 26004 6140
rect 31662 6128 31668 6140
rect 31720 6128 31726 6180
rect 32493 6171 32551 6177
rect 32493 6168 32505 6171
rect 32140 6140 32505 6168
rect 23952 6072 26004 6100
rect 26510 6060 26516 6112
rect 26568 6100 26574 6112
rect 27617 6103 27675 6109
rect 27617 6100 27629 6103
rect 26568 6072 27629 6100
rect 26568 6060 26574 6072
rect 27617 6069 27629 6072
rect 27663 6069 27675 6103
rect 27617 6063 27675 6069
rect 28718 6060 28724 6112
rect 28776 6100 28782 6112
rect 31294 6100 31300 6112
rect 28776 6072 31300 6100
rect 28776 6060 28782 6072
rect 31294 6060 31300 6072
rect 31352 6100 31358 6112
rect 32140 6100 32168 6140
rect 32493 6137 32505 6140
rect 32539 6137 32551 6171
rect 32493 6131 32551 6137
rect 33321 6171 33379 6177
rect 33321 6137 33333 6171
rect 33367 6168 33379 6171
rect 33410 6168 33416 6180
rect 33367 6140 33416 6168
rect 33367 6137 33379 6140
rect 33321 6131 33379 6137
rect 33410 6128 33416 6140
rect 33468 6128 33474 6180
rect 31352 6072 32168 6100
rect 31352 6060 31358 6072
rect 33134 6060 33140 6112
rect 33192 6100 33198 6112
rect 33229 6103 33287 6109
rect 33229 6100 33241 6103
rect 33192 6072 33241 6100
rect 33192 6060 33198 6072
rect 33229 6069 33241 6072
rect 33275 6069 33287 6103
rect 33229 6063 33287 6069
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 7742 5856 7748 5908
rect 7800 5896 7806 5908
rect 9125 5899 9183 5905
rect 9125 5896 9137 5899
rect 7800 5868 9137 5896
rect 7800 5856 7806 5868
rect 9125 5865 9137 5868
rect 9171 5865 9183 5899
rect 9950 5896 9956 5908
rect 9911 5868 9956 5896
rect 9125 5859 9183 5865
rect 9950 5856 9956 5868
rect 10008 5856 10014 5908
rect 16942 5896 16948 5908
rect 11348 5868 16948 5896
rect 9217 5831 9275 5837
rect 9217 5797 9229 5831
rect 9263 5828 9275 5831
rect 9582 5828 9588 5840
rect 9263 5800 9588 5828
rect 9263 5797 9275 5800
rect 9217 5791 9275 5797
rect 9582 5788 9588 5800
rect 9640 5828 9646 5840
rect 11348 5828 11376 5868
rect 16942 5856 16948 5868
rect 17000 5856 17006 5908
rect 17770 5896 17776 5908
rect 17731 5868 17776 5896
rect 17770 5856 17776 5868
rect 17828 5856 17834 5908
rect 19426 5896 19432 5908
rect 18708 5868 19432 5896
rect 12710 5828 12716 5840
rect 9640 5800 11376 5828
rect 11440 5800 12716 5828
rect 9640 5788 9646 5800
rect 9122 5760 9128 5772
rect 9083 5732 9128 5760
rect 9122 5720 9128 5732
rect 9180 5720 9186 5772
rect 10965 5763 11023 5769
rect 10965 5760 10977 5763
rect 10152 5732 10977 5760
rect 5534 5652 5540 5704
rect 5592 5692 5598 5704
rect 10152 5701 10180 5732
rect 10965 5729 10977 5732
rect 11011 5729 11023 5763
rect 10965 5723 11023 5729
rect 9309 5695 9367 5701
rect 9309 5692 9321 5695
rect 5592 5664 9321 5692
rect 5592 5652 5598 5664
rect 9309 5661 9321 5664
rect 9355 5661 9367 5695
rect 9309 5655 9367 5661
rect 10137 5695 10195 5701
rect 10137 5661 10149 5695
rect 10183 5661 10195 5695
rect 10594 5692 10600 5704
rect 10555 5664 10600 5692
rect 10137 5655 10195 5661
rect 10594 5652 10600 5664
rect 10652 5652 10658 5704
rect 10778 5692 10784 5704
rect 10739 5664 10784 5692
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 11440 5701 11468 5800
rect 12710 5788 12716 5800
rect 12768 5788 12774 5840
rect 14642 5828 14648 5840
rect 12820 5800 14648 5828
rect 12820 5760 12848 5800
rect 14642 5788 14648 5800
rect 14700 5788 14706 5840
rect 15746 5788 15752 5840
rect 15804 5828 15810 5840
rect 17129 5831 17187 5837
rect 17129 5828 17141 5831
rect 15804 5800 17141 5828
rect 15804 5788 15810 5800
rect 17129 5797 17141 5800
rect 17175 5797 17187 5831
rect 17129 5791 17187 5797
rect 12986 5760 12992 5772
rect 11624 5732 12848 5760
rect 12947 5732 12992 5760
rect 11624 5704 11652 5732
rect 12986 5720 12992 5732
rect 13044 5720 13050 5772
rect 16114 5720 16120 5772
rect 16172 5760 16178 5772
rect 16172 5732 18000 5760
rect 16172 5720 16178 5732
rect 11425 5695 11483 5701
rect 11425 5661 11437 5695
rect 11471 5661 11483 5695
rect 11606 5692 11612 5704
rect 11567 5664 11612 5692
rect 11425 5655 11483 5661
rect 11606 5652 11612 5664
rect 11664 5652 11670 5704
rect 11793 5695 11851 5701
rect 11793 5661 11805 5695
rect 11839 5692 11851 5695
rect 11882 5692 11888 5704
rect 11839 5664 11888 5692
rect 11839 5661 11851 5664
rect 11793 5655 11851 5661
rect 11882 5652 11888 5664
rect 11940 5692 11946 5704
rect 12713 5695 12771 5701
rect 11940 5664 12434 5692
rect 11940 5652 11946 5664
rect 8941 5627 8999 5633
rect 8941 5593 8953 5627
rect 8987 5624 8999 5627
rect 10410 5624 10416 5636
rect 8987 5596 10416 5624
rect 8987 5593 8999 5596
rect 8941 5587 8999 5593
rect 10410 5584 10416 5596
rect 10468 5584 10474 5636
rect 11701 5627 11759 5633
rect 11701 5593 11713 5627
rect 11747 5593 11759 5627
rect 12406 5624 12434 5664
rect 12713 5661 12725 5695
rect 12759 5692 12771 5695
rect 12802 5692 12808 5704
rect 12759 5664 12808 5692
rect 12759 5661 12771 5664
rect 12713 5655 12771 5661
rect 12802 5652 12808 5664
rect 12860 5652 12866 5704
rect 14642 5692 14648 5704
rect 14603 5664 14648 5692
rect 14642 5652 14648 5664
rect 14700 5652 14706 5704
rect 16669 5695 16727 5701
rect 14844 5664 16620 5692
rect 14844 5624 14872 5664
rect 12406 5596 14872 5624
rect 14912 5627 14970 5633
rect 11701 5587 11759 5593
rect 14912 5593 14924 5627
rect 14958 5624 14970 5627
rect 16206 5624 16212 5636
rect 14958 5596 16212 5624
rect 14958 5593 14970 5596
rect 14912 5587 14970 5593
rect 11422 5516 11428 5568
rect 11480 5556 11486 5568
rect 11716 5556 11744 5587
rect 16206 5584 16212 5596
rect 16264 5584 16270 5636
rect 16592 5624 16620 5664
rect 16669 5661 16681 5695
rect 16715 5692 16727 5695
rect 16758 5692 16764 5704
rect 16715 5664 16764 5692
rect 16715 5661 16727 5664
rect 16669 5655 16727 5661
rect 16758 5652 16764 5664
rect 16816 5652 16822 5704
rect 17310 5692 17316 5704
rect 17271 5664 17316 5692
rect 17310 5652 17316 5664
rect 17368 5652 17374 5704
rect 17972 5701 18000 5732
rect 18708 5701 18736 5868
rect 19426 5856 19432 5868
rect 19484 5856 19490 5908
rect 20162 5856 20168 5908
rect 20220 5896 20226 5908
rect 21726 5896 21732 5908
rect 20220 5868 21732 5896
rect 20220 5856 20226 5868
rect 21726 5856 21732 5868
rect 21784 5856 21790 5908
rect 26326 5856 26332 5908
rect 26384 5896 26390 5908
rect 26697 5899 26755 5905
rect 26697 5896 26709 5899
rect 26384 5868 26709 5896
rect 26384 5856 26390 5868
rect 26697 5865 26709 5868
rect 26743 5865 26755 5899
rect 27614 5896 27620 5908
rect 26697 5859 26755 5865
rect 26804 5868 27620 5896
rect 21082 5788 21088 5840
rect 21140 5828 21146 5840
rect 24762 5828 24768 5840
rect 21140 5800 24768 5828
rect 21140 5788 21146 5800
rect 24762 5788 24768 5800
rect 24820 5788 24826 5840
rect 25130 5788 25136 5840
rect 25188 5828 25194 5840
rect 26804 5828 26832 5868
rect 27614 5856 27620 5868
rect 27672 5856 27678 5908
rect 27890 5856 27896 5908
rect 27948 5896 27954 5908
rect 28537 5899 28595 5905
rect 28537 5896 28549 5899
rect 27948 5868 28549 5896
rect 27948 5856 27954 5868
rect 28537 5865 28549 5868
rect 28583 5865 28595 5899
rect 28537 5859 28595 5865
rect 28629 5899 28687 5905
rect 28629 5865 28641 5899
rect 28675 5896 28687 5899
rect 28718 5896 28724 5908
rect 28675 5868 28724 5896
rect 28675 5865 28687 5868
rect 28629 5859 28687 5865
rect 28718 5856 28724 5868
rect 28776 5856 28782 5908
rect 28920 5868 29684 5896
rect 25188 5800 26832 5828
rect 25188 5788 25194 5800
rect 26878 5788 26884 5840
rect 26936 5788 26942 5840
rect 28810 5828 28816 5840
rect 28552 5800 28816 5828
rect 19242 5760 19248 5772
rect 19203 5732 19248 5760
rect 19242 5720 19248 5732
rect 19300 5720 19306 5772
rect 23566 5760 23572 5772
rect 22066 5732 23572 5760
rect 17957 5695 18015 5701
rect 17957 5661 17969 5695
rect 18003 5661 18015 5695
rect 17957 5655 18015 5661
rect 18693 5695 18751 5701
rect 18693 5661 18705 5695
rect 18739 5661 18751 5695
rect 18693 5655 18751 5661
rect 18874 5652 18880 5704
rect 18932 5692 18938 5704
rect 22066 5692 22094 5732
rect 23566 5720 23572 5732
rect 23624 5720 23630 5772
rect 24854 5760 24860 5772
rect 23676 5732 24860 5760
rect 18932 5664 22094 5692
rect 22373 5695 22431 5701
rect 18932 5652 18938 5664
rect 22373 5661 22385 5695
rect 22419 5692 22431 5695
rect 22554 5692 22560 5704
rect 22419 5664 22560 5692
rect 22419 5661 22431 5664
rect 22373 5655 22431 5661
rect 22554 5652 22560 5664
rect 22612 5652 22618 5704
rect 23676 5701 23704 5732
rect 24854 5720 24860 5732
rect 24912 5720 24918 5772
rect 25317 5763 25375 5769
rect 25317 5729 25329 5763
rect 25363 5760 25375 5763
rect 26896 5760 26924 5788
rect 27430 5760 27436 5772
rect 25363 5732 27436 5760
rect 25363 5729 25375 5732
rect 25317 5723 25375 5729
rect 27430 5720 27436 5732
rect 27488 5720 27494 5772
rect 28552 5769 28580 5800
rect 28810 5788 28816 5800
rect 28868 5788 28874 5840
rect 28537 5763 28595 5769
rect 28537 5729 28549 5763
rect 28583 5729 28595 5763
rect 28920 5760 28948 5868
rect 29549 5831 29607 5837
rect 29549 5797 29561 5831
rect 29595 5797 29607 5831
rect 29656 5828 29684 5868
rect 30006 5856 30012 5908
rect 30064 5896 30070 5908
rect 30837 5899 30895 5905
rect 30837 5896 30849 5899
rect 30064 5868 30849 5896
rect 30064 5856 30070 5868
rect 30837 5865 30849 5868
rect 30883 5865 30895 5899
rect 30837 5859 30895 5865
rect 34698 5856 34704 5908
rect 34756 5896 34762 5908
rect 35802 5896 35808 5908
rect 34756 5868 35808 5896
rect 34756 5856 34762 5868
rect 35802 5856 35808 5868
rect 35860 5896 35866 5908
rect 36081 5899 36139 5905
rect 36081 5896 36093 5899
rect 35860 5868 36093 5896
rect 35860 5856 35866 5868
rect 36081 5865 36093 5868
rect 36127 5865 36139 5899
rect 37918 5896 37924 5908
rect 37879 5868 37924 5896
rect 36081 5859 36139 5865
rect 37918 5856 37924 5868
rect 37976 5856 37982 5908
rect 30193 5831 30251 5837
rect 30193 5828 30205 5831
rect 29656 5800 30205 5828
rect 29549 5791 29607 5797
rect 30193 5797 30205 5800
rect 30239 5797 30251 5831
rect 30193 5791 30251 5797
rect 28537 5723 28595 5729
rect 28644 5732 28948 5760
rect 23661 5695 23719 5701
rect 23661 5661 23673 5695
rect 23707 5661 23719 5695
rect 24394 5692 24400 5704
rect 24355 5664 24400 5692
rect 23661 5655 23719 5661
rect 24394 5652 24400 5664
rect 24452 5652 24458 5704
rect 24581 5695 24639 5701
rect 24581 5661 24593 5695
rect 24627 5661 24639 5695
rect 24581 5655 24639 5661
rect 18598 5624 18604 5636
rect 16592 5596 18604 5624
rect 18598 5584 18604 5596
rect 18656 5584 18662 5636
rect 19334 5584 19340 5636
rect 19392 5624 19398 5636
rect 19490 5627 19548 5633
rect 19490 5624 19502 5627
rect 19392 5596 19502 5624
rect 19392 5584 19398 5596
rect 19490 5593 19502 5596
rect 19536 5593 19548 5627
rect 19490 5587 19548 5593
rect 20530 5584 20536 5636
rect 20588 5624 20594 5636
rect 21637 5627 21695 5633
rect 20588 5596 20760 5624
rect 20588 5584 20594 5596
rect 11974 5556 11980 5568
rect 11480 5528 11744 5556
rect 11935 5528 11980 5556
rect 11480 5516 11486 5528
rect 11974 5516 11980 5528
rect 12032 5516 12038 5568
rect 15470 5516 15476 5568
rect 15528 5556 15534 5568
rect 16025 5559 16083 5565
rect 16025 5556 16037 5559
rect 15528 5528 16037 5556
rect 15528 5516 15534 5528
rect 16025 5525 16037 5528
rect 16071 5525 16083 5559
rect 16482 5556 16488 5568
rect 16443 5528 16488 5556
rect 16025 5519 16083 5525
rect 16482 5516 16488 5528
rect 16540 5516 16546 5568
rect 18509 5559 18567 5565
rect 18509 5525 18521 5559
rect 18555 5556 18567 5559
rect 18966 5556 18972 5568
rect 18555 5528 18972 5556
rect 18555 5525 18567 5528
rect 18509 5519 18567 5525
rect 18966 5516 18972 5528
rect 19024 5516 19030 5568
rect 19978 5516 19984 5568
rect 20036 5556 20042 5568
rect 20346 5556 20352 5568
rect 20036 5528 20352 5556
rect 20036 5516 20042 5528
rect 20346 5516 20352 5528
rect 20404 5556 20410 5568
rect 20625 5559 20683 5565
rect 20625 5556 20637 5559
rect 20404 5528 20637 5556
rect 20404 5516 20410 5528
rect 20625 5525 20637 5528
rect 20671 5525 20683 5559
rect 20732 5556 20760 5596
rect 21637 5593 21649 5627
rect 21683 5624 21695 5627
rect 21818 5624 21824 5636
rect 21683 5596 21824 5624
rect 21683 5593 21695 5596
rect 21637 5587 21695 5593
rect 21818 5584 21824 5596
rect 21876 5584 21882 5636
rect 23845 5627 23903 5633
rect 23845 5593 23857 5627
rect 23891 5624 23903 5627
rect 23934 5624 23940 5636
rect 23891 5596 23940 5624
rect 23891 5593 23903 5596
rect 23845 5587 23903 5593
rect 23934 5584 23940 5596
rect 23992 5584 23998 5636
rect 24596 5624 24624 5655
rect 24762 5652 24768 5704
rect 24820 5692 24826 5704
rect 25041 5695 25099 5701
rect 25041 5692 25053 5695
rect 24820 5664 25053 5692
rect 24820 5652 24826 5664
rect 25041 5661 25053 5664
rect 25087 5661 25099 5695
rect 26326 5692 26332 5704
rect 26287 5664 26332 5692
rect 25041 5655 25099 5661
rect 26326 5652 26332 5664
rect 26384 5652 26390 5704
rect 26510 5692 26516 5704
rect 26471 5664 26516 5692
rect 26510 5652 26516 5664
rect 26568 5652 26574 5704
rect 26878 5652 26884 5704
rect 26936 5692 26942 5704
rect 27341 5695 27399 5701
rect 27341 5692 27353 5695
rect 26936 5664 27353 5692
rect 26936 5652 26942 5664
rect 27341 5661 27353 5664
rect 27387 5661 27399 5695
rect 27341 5655 27399 5661
rect 27706 5652 27712 5704
rect 27764 5692 27770 5704
rect 28644 5692 28672 5732
rect 27764 5664 28672 5692
rect 28721 5695 28779 5701
rect 27764 5652 27770 5664
rect 28721 5661 28733 5695
rect 28767 5692 28779 5695
rect 29564 5692 29592 5791
rect 30558 5788 30564 5840
rect 30616 5828 30622 5840
rect 31481 5831 31539 5837
rect 31481 5828 31493 5831
rect 30616 5800 31493 5828
rect 30616 5788 30622 5800
rect 31481 5797 31493 5800
rect 31527 5797 31539 5831
rect 31481 5791 31539 5797
rect 28767 5664 29592 5692
rect 29733 5695 29791 5701
rect 28767 5661 28779 5664
rect 28721 5655 28779 5661
rect 29733 5661 29745 5695
rect 29779 5661 29791 5695
rect 29733 5655 29791 5661
rect 26418 5624 26424 5636
rect 24320 5596 26424 5624
rect 22278 5556 22284 5568
rect 20732 5528 22284 5556
rect 20625 5519 20683 5525
rect 22278 5516 22284 5528
rect 22336 5516 22342 5568
rect 22465 5559 22523 5565
rect 22465 5525 22477 5559
rect 22511 5556 22523 5559
rect 24320 5556 24348 5596
rect 26418 5584 26424 5596
rect 26476 5584 26482 5636
rect 28353 5627 28411 5633
rect 28353 5624 28365 5627
rect 26712 5596 28365 5624
rect 24486 5556 24492 5568
rect 22511 5528 24348 5556
rect 24447 5528 24492 5556
rect 22511 5525 22523 5528
rect 22465 5519 22523 5525
rect 24486 5516 24492 5528
rect 24544 5516 24550 5568
rect 26234 5516 26240 5568
rect 26292 5556 26298 5568
rect 26712 5556 26740 5596
rect 28353 5593 28365 5596
rect 28399 5593 28411 5627
rect 28353 5587 28411 5593
rect 26292 5528 26740 5556
rect 26292 5516 26298 5528
rect 26786 5516 26792 5568
rect 26844 5556 26850 5568
rect 27157 5559 27215 5565
rect 27157 5556 27169 5559
rect 26844 5528 27169 5556
rect 26844 5516 26850 5528
rect 27157 5525 27169 5528
rect 27203 5525 27215 5559
rect 28368 5556 28396 5587
rect 29086 5584 29092 5636
rect 29144 5624 29150 5636
rect 29748 5624 29776 5655
rect 29914 5652 29920 5704
rect 29972 5692 29978 5704
rect 30377 5695 30435 5701
rect 30377 5692 30389 5695
rect 29972 5664 30389 5692
rect 29972 5652 29978 5664
rect 30377 5661 30389 5664
rect 30423 5661 30435 5695
rect 31021 5695 31079 5701
rect 31021 5692 31033 5695
rect 30377 5655 30435 5661
rect 30484 5664 31033 5692
rect 30484 5624 30512 5664
rect 31021 5661 31033 5664
rect 31067 5661 31079 5695
rect 31021 5655 31079 5661
rect 31665 5695 31723 5701
rect 31665 5661 31677 5695
rect 31711 5661 31723 5695
rect 32306 5692 32312 5704
rect 32267 5664 32312 5692
rect 31665 5655 31723 5661
rect 29144 5596 29776 5624
rect 29840 5596 30512 5624
rect 29144 5584 29150 5596
rect 29546 5556 29552 5568
rect 28368 5528 29552 5556
rect 27157 5519 27215 5525
rect 29546 5516 29552 5528
rect 29604 5516 29610 5568
rect 29730 5516 29736 5568
rect 29788 5556 29794 5568
rect 29840 5556 29868 5596
rect 30926 5584 30932 5636
rect 30984 5624 30990 5636
rect 31680 5624 31708 5655
rect 32306 5652 32312 5664
rect 32364 5652 32370 5704
rect 34701 5695 34759 5701
rect 34701 5692 34713 5695
rect 33612 5664 34713 5692
rect 30984 5596 31708 5624
rect 30984 5584 30990 5596
rect 29788 5528 29868 5556
rect 29788 5516 29794 5528
rect 30374 5516 30380 5568
rect 30432 5556 30438 5568
rect 31110 5556 31116 5568
rect 30432 5528 31116 5556
rect 30432 5516 30438 5528
rect 31110 5516 31116 5528
rect 31168 5516 31174 5568
rect 32122 5516 32128 5568
rect 32180 5556 32186 5568
rect 33612 5565 33640 5664
rect 34701 5661 34713 5664
rect 34747 5661 34759 5695
rect 34701 5655 34759 5661
rect 38105 5695 38163 5701
rect 38105 5661 38117 5695
rect 38151 5692 38163 5695
rect 39022 5692 39028 5704
rect 38151 5664 39028 5692
rect 38151 5661 38163 5664
rect 38105 5655 38163 5661
rect 39022 5652 39028 5664
rect 39080 5652 39086 5704
rect 34514 5584 34520 5636
rect 34572 5624 34578 5636
rect 34946 5627 35004 5633
rect 34946 5624 34958 5627
rect 34572 5596 34958 5624
rect 34572 5584 34578 5596
rect 34946 5593 34958 5596
rect 34992 5593 35004 5627
rect 34946 5587 35004 5593
rect 33597 5559 33655 5565
rect 33597 5556 33609 5559
rect 32180 5528 33609 5556
rect 32180 5516 32186 5528
rect 33597 5525 33609 5528
rect 33643 5525 33655 5559
rect 33597 5519 33655 5525
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 9490 5352 9496 5364
rect 9451 5324 9496 5352
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 10502 5312 10508 5364
rect 10560 5352 10566 5364
rect 10597 5355 10655 5361
rect 10597 5352 10609 5355
rect 10560 5324 10609 5352
rect 10560 5312 10566 5324
rect 10597 5321 10609 5324
rect 10643 5321 10655 5355
rect 11698 5352 11704 5364
rect 11659 5324 11704 5352
rect 10597 5315 10655 5321
rect 11698 5312 11704 5324
rect 11756 5312 11762 5364
rect 18693 5355 18751 5361
rect 18693 5321 18705 5355
rect 18739 5352 18751 5355
rect 18782 5352 18788 5364
rect 18739 5324 18788 5352
rect 18739 5321 18751 5324
rect 18693 5315 18751 5321
rect 18782 5312 18788 5324
rect 18840 5312 18846 5364
rect 20070 5312 20076 5364
rect 20128 5352 20134 5364
rect 22186 5352 22192 5364
rect 20128 5324 22192 5352
rect 20128 5312 20134 5324
rect 22186 5312 22192 5324
rect 22244 5312 22250 5364
rect 26421 5355 26479 5361
rect 26421 5321 26433 5355
rect 26467 5352 26479 5355
rect 31573 5355 31631 5361
rect 26467 5324 27108 5352
rect 26467 5321 26479 5324
rect 26421 5315 26479 5321
rect 8754 5244 8760 5296
rect 8812 5284 8818 5296
rect 14369 5287 14427 5293
rect 14369 5284 14381 5287
rect 8812 5256 14381 5284
rect 8812 5244 8818 5256
rect 14369 5253 14381 5256
rect 14415 5253 14427 5287
rect 14369 5247 14427 5253
rect 20162 5244 20168 5296
rect 20220 5284 20226 5296
rect 20993 5287 21051 5293
rect 20220 5256 20484 5284
rect 20220 5244 20226 5256
rect 9677 5219 9735 5225
rect 9677 5185 9689 5219
rect 9723 5216 9735 5219
rect 10226 5216 10232 5228
rect 9723 5188 10232 5216
rect 9723 5185 9735 5188
rect 9677 5179 9735 5185
rect 10226 5176 10232 5188
rect 10284 5176 10290 5228
rect 10502 5176 10508 5228
rect 10560 5216 10566 5228
rect 10781 5219 10839 5225
rect 10781 5216 10793 5219
rect 10560 5188 10793 5216
rect 10560 5176 10566 5188
rect 10781 5185 10793 5188
rect 10827 5185 10839 5219
rect 10781 5179 10839 5185
rect 11606 5176 11612 5228
rect 11664 5216 11670 5228
rect 11885 5219 11943 5225
rect 11885 5216 11897 5219
rect 11664 5188 11897 5216
rect 11664 5176 11670 5188
rect 11885 5185 11897 5188
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 12796 5219 12854 5225
rect 12796 5185 12808 5219
rect 12842 5216 12854 5219
rect 13998 5216 14004 5228
rect 12842 5188 14004 5216
rect 12842 5185 12854 5188
rect 12796 5179 12854 5185
rect 13998 5176 14004 5188
rect 14056 5176 14062 5228
rect 17218 5216 17224 5228
rect 17179 5188 17224 5216
rect 17218 5176 17224 5188
rect 17276 5176 17282 5228
rect 17405 5219 17463 5225
rect 17405 5185 17417 5219
rect 17451 5185 17463 5219
rect 17405 5179 17463 5185
rect 12434 5108 12440 5160
rect 12492 5148 12498 5160
rect 12529 5151 12587 5157
rect 12529 5148 12541 5151
rect 12492 5120 12541 5148
rect 12492 5108 12498 5120
rect 12529 5117 12541 5120
rect 12575 5117 12587 5151
rect 12529 5111 12587 5117
rect 12544 5012 12572 5111
rect 13538 5108 13544 5160
rect 13596 5148 13602 5160
rect 14642 5148 14648 5160
rect 13596 5120 14648 5148
rect 13596 5108 13602 5120
rect 14642 5108 14648 5120
rect 14700 5148 14706 5160
rect 16117 5151 16175 5157
rect 16117 5148 16129 5151
rect 14700 5120 16129 5148
rect 14700 5108 14706 5120
rect 16117 5117 16129 5120
rect 16163 5148 16175 5151
rect 16850 5148 16856 5160
rect 16163 5120 16856 5148
rect 16163 5117 16175 5120
rect 16117 5111 16175 5117
rect 16850 5108 16856 5120
rect 16908 5108 16914 5160
rect 16298 5040 16304 5092
rect 16356 5080 16362 5092
rect 17420 5080 17448 5179
rect 17954 5176 17960 5228
rect 18012 5216 18018 5228
rect 18233 5219 18291 5225
rect 18233 5216 18245 5219
rect 18012 5188 18245 5216
rect 18012 5176 18018 5188
rect 18233 5185 18245 5188
rect 18279 5185 18291 5219
rect 18233 5179 18291 5185
rect 18414 5176 18420 5228
rect 18472 5216 18478 5228
rect 18877 5219 18935 5225
rect 18877 5216 18889 5219
rect 18472 5188 18889 5216
rect 18472 5176 18478 5188
rect 18877 5185 18889 5188
rect 18923 5185 18935 5219
rect 18877 5179 18935 5185
rect 19242 5176 19248 5228
rect 19300 5216 19306 5228
rect 20456 5225 20484 5256
rect 20993 5253 21005 5287
rect 21039 5284 21051 5287
rect 22554 5284 22560 5296
rect 21039 5256 22560 5284
rect 21039 5253 21051 5256
rect 20993 5247 21051 5253
rect 22554 5244 22560 5256
rect 22612 5244 22618 5296
rect 25038 5284 25044 5296
rect 23400 5256 25044 5284
rect 19407 5219 19465 5225
rect 19407 5216 19419 5219
rect 19300 5188 19419 5216
rect 19300 5176 19306 5188
rect 19407 5185 19419 5188
rect 19453 5185 19465 5219
rect 19407 5179 19465 5185
rect 19705 5219 19763 5225
rect 19705 5185 19717 5219
rect 19751 5216 19763 5219
rect 20441 5219 20499 5225
rect 19751 5188 20300 5216
rect 19751 5185 19763 5188
rect 19705 5179 19763 5185
rect 19521 5151 19579 5157
rect 19521 5117 19533 5151
rect 19567 5148 19579 5151
rect 19978 5148 19984 5160
rect 19567 5120 19984 5148
rect 19567 5117 19579 5120
rect 19521 5111 19579 5117
rect 19978 5108 19984 5120
rect 20036 5108 20042 5160
rect 16356 5052 17448 5080
rect 16356 5040 16362 5052
rect 17770 5040 17776 5092
rect 17828 5080 17834 5092
rect 19337 5083 19395 5089
rect 19337 5080 19349 5083
rect 17828 5052 19349 5080
rect 17828 5040 17834 5052
rect 19337 5049 19349 5052
rect 19383 5080 19395 5083
rect 19702 5080 19708 5092
rect 19383 5052 19708 5080
rect 19383 5049 19395 5052
rect 19337 5043 19395 5049
rect 19702 5040 19708 5052
rect 19760 5040 19766 5092
rect 20272 5089 20300 5188
rect 20441 5185 20453 5219
rect 20487 5185 20499 5219
rect 20441 5179 20499 5185
rect 21266 5176 21272 5228
rect 21324 5216 21330 5228
rect 22005 5219 22063 5225
rect 22005 5216 22017 5219
rect 21324 5188 22017 5216
rect 21324 5176 21330 5188
rect 22005 5185 22017 5188
rect 22051 5185 22063 5219
rect 22005 5179 22063 5185
rect 22741 5219 22799 5225
rect 22741 5185 22753 5219
rect 22787 5216 22799 5219
rect 23198 5216 23204 5228
rect 22787 5188 23204 5216
rect 22787 5185 22799 5188
rect 22741 5179 22799 5185
rect 23198 5176 23204 5188
rect 23256 5176 23262 5228
rect 23400 5225 23428 5256
rect 25038 5244 25044 5256
rect 25096 5244 25102 5296
rect 27080 5284 27108 5324
rect 27540 5324 30788 5352
rect 27218 5287 27276 5293
rect 27218 5284 27230 5287
rect 27080 5256 27230 5284
rect 27218 5253 27230 5256
rect 27264 5253 27276 5287
rect 27218 5247 27276 5253
rect 27540 5228 27568 5324
rect 29638 5284 29644 5296
rect 28828 5256 29644 5284
rect 23385 5219 23443 5225
rect 23385 5185 23397 5219
rect 23431 5185 23443 5219
rect 23385 5179 23443 5185
rect 23652 5219 23710 5225
rect 23652 5185 23664 5219
rect 23698 5216 23710 5219
rect 24486 5216 24492 5228
rect 23698 5188 24492 5216
rect 23698 5185 23710 5188
rect 23652 5179 23710 5185
rect 24486 5176 24492 5188
rect 24544 5176 24550 5228
rect 25317 5219 25375 5225
rect 25317 5185 25329 5219
rect 25363 5185 25375 5219
rect 26234 5216 26240 5228
rect 26195 5188 26240 5216
rect 25317 5179 25375 5185
rect 25332 5148 25360 5179
rect 26234 5176 26240 5188
rect 26292 5176 26298 5228
rect 26418 5216 26424 5228
rect 26379 5188 26424 5216
rect 26418 5176 26424 5188
rect 26476 5216 26482 5228
rect 27522 5216 27528 5228
rect 26476 5188 27528 5216
rect 26476 5176 26482 5188
rect 27522 5176 27528 5188
rect 27580 5176 27586 5228
rect 28828 5225 28856 5256
rect 29638 5244 29644 5256
rect 29696 5244 29702 5296
rect 28813 5219 28871 5225
rect 28813 5185 28825 5219
rect 28859 5185 28871 5219
rect 29069 5219 29127 5225
rect 29069 5216 29081 5219
rect 28813 5179 28871 5185
rect 28920 5188 29081 5216
rect 26970 5148 26976 5160
rect 24504 5120 25360 5148
rect 26931 5120 26976 5148
rect 20257 5083 20315 5089
rect 20257 5049 20269 5083
rect 20303 5049 20315 5083
rect 20257 5043 20315 5049
rect 20990 5040 20996 5092
rect 21048 5080 21054 5092
rect 21821 5083 21879 5089
rect 21821 5080 21833 5083
rect 21048 5052 21833 5080
rect 21048 5040 21054 5052
rect 21821 5049 21833 5052
rect 21867 5049 21879 5083
rect 21821 5043 21879 5049
rect 13538 5012 13544 5024
rect 12544 4984 13544 5012
rect 13538 4972 13544 4984
rect 13596 4972 13602 5024
rect 13909 5015 13967 5021
rect 13909 4981 13921 5015
rect 13955 5012 13967 5015
rect 14274 5012 14280 5024
rect 13955 4984 14280 5012
rect 13955 4981 13967 4984
rect 13909 4975 13967 4981
rect 14274 4972 14280 4984
rect 14332 4972 14338 5024
rect 17310 5012 17316 5024
rect 17271 4984 17316 5012
rect 17310 4972 17316 4984
rect 17368 4972 17374 5024
rect 18046 5012 18052 5024
rect 18007 4984 18052 5012
rect 18046 4972 18052 4984
rect 18104 4972 18110 5024
rect 18966 4972 18972 5024
rect 19024 5012 19030 5024
rect 19613 5015 19671 5021
rect 19613 5012 19625 5015
rect 19024 4984 19625 5012
rect 19024 4972 19030 4984
rect 19613 4981 19625 4984
rect 19659 4981 19671 5015
rect 19613 4975 19671 4981
rect 20898 4972 20904 5024
rect 20956 5012 20962 5024
rect 21085 5015 21143 5021
rect 21085 5012 21097 5015
rect 20956 4984 21097 5012
rect 20956 4972 20962 4984
rect 21085 4981 21097 4984
rect 21131 4981 21143 5015
rect 21085 4975 21143 4981
rect 22002 4972 22008 5024
rect 22060 5012 22066 5024
rect 22833 5015 22891 5021
rect 22833 5012 22845 5015
rect 22060 4984 22845 5012
rect 22060 4972 22066 4984
rect 22833 4981 22845 4984
rect 22879 4981 22891 5015
rect 22833 4975 22891 4981
rect 23198 4972 23204 5024
rect 23256 5012 23262 5024
rect 24504 5012 24532 5120
rect 26970 5108 26976 5120
rect 27028 5108 27034 5160
rect 27982 5108 27988 5160
rect 28040 5148 28046 5160
rect 28920 5148 28948 5188
rect 29069 5185 29081 5188
rect 29115 5185 29127 5219
rect 29069 5179 29127 5185
rect 30466 5176 30472 5228
rect 30524 5216 30530 5228
rect 30653 5219 30711 5225
rect 30653 5216 30665 5219
rect 30524 5188 30665 5216
rect 30524 5176 30530 5188
rect 30653 5185 30665 5188
rect 30699 5185 30711 5219
rect 30760 5216 30788 5324
rect 31573 5321 31585 5355
rect 31619 5352 31631 5355
rect 34425 5355 34483 5361
rect 31619 5324 32076 5352
rect 31619 5321 31631 5324
rect 31573 5315 31631 5321
rect 31938 5284 31944 5296
rect 31404 5256 31944 5284
rect 31404 5225 31432 5256
rect 31938 5244 31944 5256
rect 31996 5244 32002 5296
rect 32048 5284 32076 5324
rect 34425 5321 34437 5355
rect 34471 5352 34483 5355
rect 34514 5352 34520 5364
rect 34471 5324 34520 5352
rect 34471 5321 34483 5324
rect 34425 5315 34483 5321
rect 34514 5312 34520 5324
rect 34572 5312 34578 5364
rect 32370 5287 32428 5293
rect 32370 5284 32382 5287
rect 32048 5256 32382 5284
rect 32370 5253 32382 5256
rect 32416 5253 32428 5287
rect 32370 5247 32428 5253
rect 30837 5219 30895 5225
rect 30837 5216 30849 5219
rect 30760 5188 30849 5216
rect 30653 5179 30711 5185
rect 30837 5185 30849 5188
rect 30883 5185 30895 5219
rect 30837 5179 30895 5185
rect 31389 5219 31447 5225
rect 31389 5185 31401 5219
rect 31435 5185 31447 5219
rect 31389 5179 31447 5185
rect 31573 5219 31631 5225
rect 31573 5185 31585 5219
rect 31619 5185 31631 5219
rect 31573 5179 31631 5185
rect 28040 5120 28948 5148
rect 30852 5148 30880 5179
rect 31588 5148 31616 5179
rect 31846 5176 31852 5228
rect 31904 5216 31910 5228
rect 34606 5216 34612 5228
rect 31904 5188 33456 5216
rect 34567 5188 34612 5216
rect 31904 5176 31910 5188
rect 32122 5148 32128 5160
rect 30852 5120 31616 5148
rect 32035 5120 32128 5148
rect 28040 5108 28046 5120
rect 32122 5108 32128 5120
rect 32180 5108 32186 5160
rect 31570 5040 31576 5092
rect 31628 5080 31634 5092
rect 32140 5080 32168 5108
rect 31628 5052 32168 5080
rect 33428 5080 33456 5188
rect 34606 5176 34612 5188
rect 34664 5176 34670 5228
rect 35253 5219 35311 5225
rect 35253 5185 35265 5219
rect 35299 5216 35311 5219
rect 35342 5216 35348 5228
rect 35299 5188 35348 5216
rect 35299 5185 35311 5188
rect 35253 5179 35311 5185
rect 35342 5176 35348 5188
rect 35400 5176 35406 5228
rect 37826 5216 37832 5228
rect 37787 5188 37832 5216
rect 37826 5176 37832 5188
rect 37884 5176 37890 5228
rect 35069 5083 35127 5089
rect 35069 5080 35081 5083
rect 33428 5052 35081 5080
rect 31628 5040 31634 5052
rect 35069 5049 35081 5052
rect 35115 5049 35127 5083
rect 35069 5043 35127 5049
rect 23256 4984 24532 5012
rect 23256 4972 23262 4984
rect 24578 4972 24584 5024
rect 24636 5012 24642 5024
rect 24765 5015 24823 5021
rect 24765 5012 24777 5015
rect 24636 4984 24777 5012
rect 24636 4972 24642 4984
rect 24765 4981 24777 4984
rect 24811 4981 24823 5015
rect 25406 5012 25412 5024
rect 25319 4984 25412 5012
rect 24765 4975 24823 4981
rect 25406 4972 25412 4984
rect 25464 5012 25470 5024
rect 27614 5012 27620 5024
rect 25464 4984 27620 5012
rect 25464 4972 25470 4984
rect 27614 4972 27620 4984
rect 27672 4972 27678 5024
rect 28350 5012 28356 5024
rect 28311 4984 28356 5012
rect 28350 4972 28356 4984
rect 28408 4972 28414 5024
rect 28810 4972 28816 5024
rect 28868 5012 28874 5024
rect 30193 5015 30251 5021
rect 30193 5012 30205 5015
rect 28868 4984 30205 5012
rect 28868 4972 28874 4984
rect 30193 4981 30205 4984
rect 30239 4981 30251 5015
rect 30742 5012 30748 5024
rect 30703 4984 30748 5012
rect 30193 4975 30251 4981
rect 30742 4972 30748 4984
rect 30800 4972 30806 5024
rect 32398 4972 32404 5024
rect 32456 5012 32462 5024
rect 33505 5015 33563 5021
rect 33505 5012 33517 5015
rect 32456 4984 33517 5012
rect 32456 4972 32462 4984
rect 33505 4981 33517 4984
rect 33551 4981 33563 5015
rect 33505 4975 33563 4981
rect 38013 5015 38071 5021
rect 38013 4981 38025 5015
rect 38059 5012 38071 5015
rect 39758 5012 39764 5024
rect 38059 4984 39764 5012
rect 38059 4981 38071 4984
rect 38013 4975 38071 4981
rect 39758 4972 39764 4984
rect 39816 4972 39822 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 10410 4768 10416 4820
rect 10468 4808 10474 4820
rect 10468 4780 12434 4808
rect 10468 4768 10474 4780
rect 10229 4743 10287 4749
rect 10229 4709 10241 4743
rect 10275 4740 10287 4743
rect 11790 4740 11796 4752
rect 10275 4712 11796 4740
rect 10275 4709 10287 4712
rect 10229 4703 10287 4709
rect 11790 4700 11796 4712
rect 11848 4700 11854 4752
rect 12406 4740 12434 4780
rect 13906 4768 13912 4820
rect 13964 4808 13970 4820
rect 14277 4811 14335 4817
rect 14277 4808 14289 4811
rect 13964 4780 14289 4808
rect 13964 4768 13970 4780
rect 14277 4777 14289 4780
rect 14323 4777 14335 4811
rect 14277 4771 14335 4777
rect 14369 4811 14427 4817
rect 14369 4777 14381 4811
rect 14415 4808 14427 4811
rect 15565 4811 15623 4817
rect 15565 4808 15577 4811
rect 14415 4780 15577 4808
rect 14415 4777 14427 4780
rect 14369 4771 14427 4777
rect 15565 4777 15577 4780
rect 15611 4808 15623 4811
rect 17586 4808 17592 4820
rect 15611 4780 17592 4808
rect 15611 4777 15623 4780
rect 15565 4771 15623 4777
rect 17586 4768 17592 4780
rect 17644 4808 17650 4820
rect 18966 4808 18972 4820
rect 17644 4780 18972 4808
rect 17644 4768 17650 4780
rect 18966 4768 18972 4780
rect 19024 4768 19030 4820
rect 19334 4808 19340 4820
rect 19295 4780 19340 4808
rect 19334 4768 19340 4780
rect 19392 4768 19398 4820
rect 22002 4768 22008 4820
rect 22060 4808 22066 4820
rect 22060 4780 22105 4808
rect 22060 4768 22066 4780
rect 24394 4768 24400 4820
rect 24452 4808 24458 4820
rect 24581 4811 24639 4817
rect 24581 4808 24593 4811
rect 24452 4780 24593 4808
rect 24452 4768 24458 4780
rect 24581 4777 24593 4780
rect 24627 4777 24639 4811
rect 24581 4771 24639 4777
rect 24673 4811 24731 4817
rect 24673 4777 24685 4811
rect 24719 4808 24731 4811
rect 25406 4808 25412 4820
rect 24719 4780 25412 4808
rect 24719 4777 24731 4780
rect 24673 4771 24731 4777
rect 25406 4768 25412 4780
rect 25464 4768 25470 4820
rect 26234 4768 26240 4820
rect 26292 4808 26298 4820
rect 26605 4811 26663 4817
rect 26605 4808 26617 4811
rect 26292 4780 26617 4808
rect 26292 4768 26298 4780
rect 26605 4777 26617 4780
rect 26651 4777 26663 4811
rect 26605 4771 26663 4777
rect 26697 4811 26755 4817
rect 26697 4777 26709 4811
rect 26743 4808 26755 4811
rect 27614 4808 27620 4820
rect 26743 4780 27620 4808
rect 26743 4777 26755 4780
rect 26697 4771 26755 4777
rect 27614 4768 27620 4780
rect 27672 4808 27678 4820
rect 27982 4808 27988 4820
rect 27672 4780 27844 4808
rect 27943 4780 27988 4808
rect 27672 4768 27678 4780
rect 14093 4743 14151 4749
rect 14093 4740 14105 4743
rect 12406 4712 14105 4740
rect 14093 4709 14105 4712
rect 14139 4740 14151 4743
rect 14182 4740 14188 4752
rect 14139 4712 14188 4740
rect 14139 4709 14151 4712
rect 14093 4703 14151 4709
rect 14182 4700 14188 4712
rect 14240 4700 14246 4752
rect 15359 4743 15417 4749
rect 15359 4709 15371 4743
rect 15405 4740 15417 4743
rect 18984 4740 19012 4768
rect 20806 4740 20812 4752
rect 15405 4712 16160 4740
rect 18984 4712 20812 4740
rect 15405 4709 15417 4712
rect 15359 4703 15417 4709
rect 14274 4672 14280 4684
rect 14235 4644 14280 4672
rect 14274 4632 14280 4644
rect 14332 4632 14338 4684
rect 15470 4672 15476 4684
rect 15431 4644 15476 4672
rect 15470 4632 15476 4644
rect 15528 4632 15534 4684
rect 15580 4644 15792 4672
rect 9033 4607 9091 4613
rect 9033 4573 9045 4607
rect 9079 4573 9091 4607
rect 9033 4567 9091 4573
rect 9048 4536 9076 4567
rect 9122 4564 9128 4616
rect 9180 4604 9186 4616
rect 9217 4607 9275 4613
rect 9217 4604 9229 4607
rect 9180 4576 9229 4604
rect 9180 4564 9186 4576
rect 9217 4573 9229 4576
rect 9263 4604 9275 4607
rect 9306 4604 9312 4616
rect 9263 4576 9312 4604
rect 9263 4573 9275 4576
rect 9217 4567 9275 4573
rect 9306 4564 9312 4576
rect 9364 4564 9370 4616
rect 10134 4564 10140 4616
rect 10192 4604 10198 4616
rect 10413 4607 10471 4613
rect 10413 4604 10425 4607
rect 10192 4576 10425 4604
rect 10192 4564 10198 4576
rect 10413 4573 10425 4576
rect 10459 4573 10471 4607
rect 10413 4567 10471 4573
rect 11238 4564 11244 4616
rect 11296 4604 11302 4616
rect 11517 4607 11575 4613
rect 11517 4604 11529 4607
rect 11296 4576 11529 4604
rect 11296 4564 11302 4576
rect 11517 4573 11529 4576
rect 11563 4573 11575 4607
rect 11517 4567 11575 4573
rect 12253 4607 12311 4613
rect 12253 4573 12265 4607
rect 12299 4604 12311 4607
rect 12434 4604 12440 4616
rect 12299 4576 12440 4604
rect 12299 4573 12311 4576
rect 12253 4567 12311 4573
rect 12434 4564 12440 4576
rect 12492 4564 12498 4616
rect 12618 4564 12624 4616
rect 12676 4604 12682 4616
rect 12897 4607 12955 4613
rect 12897 4604 12909 4607
rect 12676 4576 12909 4604
rect 12676 4564 12682 4576
rect 12897 4573 12909 4576
rect 12943 4573 12955 4607
rect 12897 4567 12955 4573
rect 13541 4607 13599 4613
rect 13541 4573 13553 4607
rect 13587 4604 13599 4607
rect 14182 4604 14188 4616
rect 13587 4576 14188 4604
rect 13587 4573 13599 4576
rect 13541 4567 13599 4573
rect 14182 4564 14188 4576
rect 14240 4564 14246 4616
rect 14461 4607 14519 4613
rect 14461 4573 14473 4607
rect 14507 4604 14519 4607
rect 15580 4604 15608 4644
rect 14507 4576 15608 4604
rect 15657 4607 15715 4613
rect 14507 4573 14519 4576
rect 14461 4567 14519 4573
rect 15657 4573 15669 4607
rect 15703 4573 15715 4607
rect 15657 4567 15715 4573
rect 10594 4536 10600 4548
rect 9048 4508 10600 4536
rect 10594 4496 10600 4508
rect 10652 4496 10658 4548
rect 15286 4536 15292 4548
rect 15247 4508 15292 4536
rect 15286 4496 15292 4508
rect 15344 4496 15350 4548
rect 9122 4468 9128 4480
rect 9083 4440 9128 4468
rect 9122 4428 9128 4440
rect 9180 4428 9186 4480
rect 11330 4468 11336 4480
rect 11291 4440 11336 4468
rect 11330 4428 11336 4440
rect 11388 4428 11394 4480
rect 12066 4468 12072 4480
rect 12027 4440 12072 4468
rect 12066 4428 12072 4440
rect 12124 4428 12130 4480
rect 12713 4471 12771 4477
rect 12713 4437 12725 4471
rect 12759 4468 12771 4471
rect 12802 4468 12808 4480
rect 12759 4440 12808 4468
rect 12759 4437 12771 4440
rect 12713 4431 12771 4437
rect 12802 4428 12808 4440
rect 12860 4428 12866 4480
rect 13354 4468 13360 4480
rect 13315 4440 13360 4468
rect 13354 4428 13360 4440
rect 13412 4428 13418 4480
rect 15672 4468 15700 4567
rect 15764 4536 15792 4644
rect 16132 4613 16160 4712
rect 20806 4700 20812 4712
rect 20864 4700 20870 4752
rect 27249 4743 27307 4749
rect 27249 4740 27261 4743
rect 24872 4712 27261 4740
rect 16206 4632 16212 4684
rect 16264 4672 16270 4684
rect 20898 4672 20904 4684
rect 16264 4644 16309 4672
rect 19444 4644 20904 4672
rect 16264 4632 16270 4644
rect 16117 4607 16175 4613
rect 16117 4573 16129 4607
rect 16163 4573 16175 4607
rect 16298 4604 16304 4616
rect 16259 4576 16304 4604
rect 16117 4567 16175 4573
rect 16298 4564 16304 4576
rect 16356 4604 16362 4616
rect 16850 4604 16856 4616
rect 16356 4576 16712 4604
rect 16763 4576 16856 4604
rect 16356 4564 16362 4576
rect 16482 4536 16488 4548
rect 15764 4508 16488 4536
rect 16482 4496 16488 4508
rect 16540 4496 16546 4548
rect 16684 4536 16712 4576
rect 16850 4564 16856 4576
rect 16908 4604 16914 4616
rect 17862 4604 17868 4616
rect 16908 4576 17868 4604
rect 16908 4564 16914 4576
rect 17862 4564 17868 4576
rect 17920 4564 17926 4616
rect 19242 4604 19248 4616
rect 19203 4576 19248 4604
rect 19242 4564 19248 4576
rect 19300 4564 19306 4616
rect 19444 4613 19472 4644
rect 20898 4632 20904 4644
rect 20956 4672 20962 4684
rect 21726 4672 21732 4684
rect 20956 4644 21220 4672
rect 21687 4644 21732 4672
rect 20956 4632 20962 4644
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4573 19487 4607
rect 20070 4604 20076 4616
rect 20031 4576 20076 4604
rect 19429 4567 19487 4573
rect 17120 4539 17178 4545
rect 16684 4508 17080 4536
rect 16942 4468 16948 4480
rect 15672 4440 16948 4468
rect 16942 4428 16948 4440
rect 17000 4428 17006 4480
rect 17052 4468 17080 4508
rect 17120 4505 17132 4539
rect 17166 4536 17178 4539
rect 17310 4536 17316 4548
rect 17166 4508 17316 4536
rect 17166 4505 17178 4508
rect 17120 4499 17178 4505
rect 17310 4496 17316 4508
rect 17368 4496 17374 4548
rect 19444 4536 19472 4567
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 21085 4607 21143 4613
rect 21085 4573 21097 4607
rect 21131 4573 21143 4607
rect 21085 4567 21143 4573
rect 21192 4600 21220 4644
rect 21726 4632 21732 4644
rect 21784 4632 21790 4684
rect 21867 4675 21925 4681
rect 21867 4641 21879 4675
rect 21913 4641 21925 4675
rect 21867 4635 21925 4641
rect 21269 4607 21327 4613
rect 21269 4600 21281 4607
rect 21192 4573 21281 4600
rect 21315 4573 21327 4607
rect 21192 4572 21327 4573
rect 21882 4600 21910 4635
rect 22186 4632 22192 4684
rect 22244 4672 22250 4684
rect 22244 4644 22600 4672
rect 22244 4632 22250 4644
rect 22002 4600 22008 4616
rect 21882 4572 22008 4600
rect 21269 4567 21327 4572
rect 18064 4508 19472 4536
rect 21100 4536 21128 4567
rect 22002 4564 22008 4572
rect 22060 4564 22066 4616
rect 22097 4607 22155 4613
rect 22097 4573 22109 4607
rect 22143 4604 22155 4607
rect 22462 4604 22468 4616
rect 22143 4576 22468 4604
rect 22143 4573 22155 4576
rect 22097 4567 22155 4573
rect 22462 4564 22468 4576
rect 22520 4564 22526 4616
rect 22572 4613 22600 4644
rect 23934 4632 23940 4684
rect 23992 4672 23998 4684
rect 24397 4675 24455 4681
rect 24397 4672 24409 4675
rect 23992 4644 24409 4672
rect 23992 4632 23998 4644
rect 24397 4641 24409 4644
rect 24443 4641 24455 4675
rect 24578 4672 24584 4684
rect 24539 4644 24584 4672
rect 24397 4635 24455 4641
rect 24578 4632 24584 4644
rect 24636 4632 24642 4684
rect 22557 4607 22615 4613
rect 22557 4573 22569 4607
rect 22603 4573 22615 4607
rect 22557 4567 22615 4573
rect 23293 4607 23351 4613
rect 23293 4573 23305 4607
rect 23339 4604 23351 4607
rect 23658 4604 23664 4616
rect 23339 4576 23664 4604
rect 23339 4573 23351 4576
rect 23293 4567 23351 4573
rect 23658 4564 23664 4576
rect 23716 4564 23722 4616
rect 24765 4607 24823 4613
rect 24765 4573 24777 4607
rect 24811 4604 24823 4607
rect 24872 4604 24900 4712
rect 27249 4709 27261 4712
rect 27295 4709 27307 4743
rect 27816 4740 27844 4780
rect 27982 4768 27988 4780
rect 28040 4768 28046 4820
rect 28810 4808 28816 4820
rect 28771 4780 28816 4808
rect 28810 4768 28816 4780
rect 28868 4768 28874 4820
rect 28902 4768 28908 4820
rect 28960 4808 28966 4820
rect 32214 4808 32220 4820
rect 28960 4780 32220 4808
rect 28960 4768 28966 4780
rect 32214 4768 32220 4780
rect 32272 4768 32278 4820
rect 32398 4808 32404 4820
rect 32359 4780 32404 4808
rect 32398 4768 32404 4780
rect 32456 4768 32462 4820
rect 33134 4768 33140 4820
rect 33192 4808 33198 4820
rect 33597 4811 33655 4817
rect 33597 4808 33609 4811
rect 33192 4780 33609 4808
rect 33192 4768 33198 4780
rect 33597 4777 33609 4780
rect 33643 4777 33655 4811
rect 35710 4808 35716 4820
rect 35671 4780 35716 4808
rect 33597 4771 33655 4777
rect 35710 4768 35716 4780
rect 35768 4768 35774 4820
rect 37182 4808 37188 4820
rect 37143 4780 37188 4808
rect 37182 4768 37188 4780
rect 37240 4768 37246 4820
rect 28718 4740 28724 4752
rect 27816 4712 28724 4740
rect 27249 4703 27307 4709
rect 28718 4700 28724 4712
rect 28776 4700 28782 4752
rect 31110 4700 31116 4752
rect 31168 4740 31174 4752
rect 32861 4743 32919 4749
rect 32861 4740 32873 4743
rect 31168 4712 32873 4740
rect 31168 4700 31174 4712
rect 32861 4709 32873 4712
rect 32907 4709 32919 4743
rect 32861 4703 32919 4709
rect 26326 4632 26332 4684
rect 26384 4672 26390 4684
rect 26421 4675 26479 4681
rect 26421 4672 26433 4675
rect 26384 4644 26433 4672
rect 26384 4632 26390 4644
rect 26421 4641 26433 4644
rect 26467 4641 26479 4675
rect 26421 4635 26479 4641
rect 26605 4675 26663 4681
rect 26605 4641 26617 4675
rect 26651 4641 26663 4675
rect 26605 4635 26663 4641
rect 25590 4604 25596 4616
rect 24811 4576 24900 4604
rect 25551 4576 25596 4604
rect 24811 4573 24823 4576
rect 24765 4567 24823 4573
rect 25590 4564 25596 4576
rect 25648 4564 25654 4616
rect 21799 4539 21857 4545
rect 21799 4536 21811 4539
rect 21100 4508 21811 4536
rect 18064 4468 18092 4508
rect 21799 4505 21811 4508
rect 21845 4505 21857 4539
rect 26620 4536 26648 4635
rect 27522 4632 27528 4684
rect 27580 4672 27586 4684
rect 32493 4675 32551 4681
rect 27580 4644 28120 4672
rect 27580 4632 27586 4644
rect 26786 4604 26792 4616
rect 26747 4576 26792 4604
rect 26786 4564 26792 4576
rect 26844 4564 26850 4616
rect 27430 4564 27436 4616
rect 27488 4604 27494 4616
rect 27890 4604 27896 4616
rect 27488 4576 27533 4604
rect 27851 4576 27896 4604
rect 27488 4564 27494 4576
rect 27890 4564 27896 4576
rect 27948 4564 27954 4616
rect 28092 4613 28120 4644
rect 32493 4641 32505 4675
rect 32539 4641 32551 4675
rect 32493 4635 32551 4641
rect 28077 4607 28135 4613
rect 28077 4573 28089 4607
rect 28123 4573 28135 4607
rect 28718 4604 28724 4616
rect 28679 4576 28724 4604
rect 28077 4567 28135 4573
rect 28718 4564 28724 4576
rect 28776 4564 28782 4616
rect 28813 4607 28871 4613
rect 28813 4573 28825 4607
rect 28859 4573 28871 4607
rect 28813 4567 28871 4573
rect 28350 4536 28356 4548
rect 26620 4508 28356 4536
rect 21799 4499 21857 4505
rect 28350 4496 28356 4508
rect 28408 4536 28414 4548
rect 28537 4539 28595 4545
rect 28537 4536 28549 4539
rect 28408 4508 28549 4536
rect 28408 4496 28414 4508
rect 28537 4505 28549 4508
rect 28583 4505 28595 4539
rect 28828 4536 28856 4567
rect 29638 4564 29644 4616
rect 29696 4604 29702 4616
rect 30101 4607 30159 4613
rect 30101 4604 30113 4607
rect 29696 4576 30113 4604
rect 29696 4564 29702 4576
rect 30101 4573 30113 4576
rect 30147 4604 30159 4607
rect 31570 4604 31576 4616
rect 30147 4576 31576 4604
rect 30147 4573 30159 4576
rect 30101 4567 30159 4573
rect 31570 4564 31576 4576
rect 31628 4564 31634 4616
rect 30368 4539 30426 4545
rect 28828 4508 30328 4536
rect 28537 4499 28595 4505
rect 18230 4468 18236 4480
rect 17052 4440 18092 4468
rect 18191 4440 18236 4468
rect 18230 4428 18236 4440
rect 18288 4428 18294 4480
rect 19889 4471 19947 4477
rect 19889 4437 19901 4471
rect 19935 4468 19947 4471
rect 19978 4468 19984 4480
rect 19935 4440 19984 4468
rect 19935 4437 19947 4440
rect 19889 4431 19947 4437
rect 19978 4428 19984 4440
rect 20036 4428 20042 4480
rect 21269 4471 21327 4477
rect 21269 4437 21281 4471
rect 21315 4468 21327 4471
rect 22186 4468 22192 4480
rect 21315 4440 22192 4468
rect 21315 4437 21327 4440
rect 21269 4431 21327 4437
rect 22186 4428 22192 4440
rect 22244 4428 22250 4480
rect 22278 4428 22284 4480
rect 22336 4468 22342 4480
rect 22741 4471 22799 4477
rect 22741 4468 22753 4471
rect 22336 4440 22753 4468
rect 22336 4428 22342 4440
rect 22741 4437 22753 4440
rect 22787 4437 22799 4471
rect 23474 4468 23480 4480
rect 23435 4440 23480 4468
rect 22741 4431 22799 4437
rect 23474 4428 23480 4440
rect 23532 4428 23538 4480
rect 25314 4428 25320 4480
rect 25372 4468 25378 4480
rect 25409 4471 25467 4477
rect 25409 4468 25421 4471
rect 25372 4440 25421 4468
rect 25372 4428 25378 4440
rect 25409 4437 25421 4440
rect 25455 4437 25467 4471
rect 25409 4431 25467 4437
rect 28997 4471 29055 4477
rect 28997 4437 29009 4471
rect 29043 4468 29055 4471
rect 29454 4468 29460 4480
rect 29043 4440 29460 4468
rect 29043 4437 29055 4440
rect 28997 4431 29055 4437
rect 29454 4428 29460 4440
rect 29512 4428 29518 4480
rect 30300 4468 30328 4508
rect 30368 4505 30380 4539
rect 30414 4536 30426 4539
rect 30742 4536 30748 4548
rect 30414 4508 30748 4536
rect 30414 4505 30426 4508
rect 30368 4499 30426 4505
rect 30742 4496 30748 4508
rect 30800 4496 30806 4548
rect 32401 4539 32459 4545
rect 32401 4536 32413 4539
rect 31726 4508 32413 4536
rect 30558 4468 30564 4480
rect 30300 4440 30564 4468
rect 30558 4428 30564 4440
rect 30616 4428 30622 4480
rect 30834 4428 30840 4480
rect 30892 4468 30898 4480
rect 31481 4471 31539 4477
rect 31481 4468 31493 4471
rect 30892 4440 31493 4468
rect 30892 4428 30898 4440
rect 31481 4437 31493 4440
rect 31527 4468 31539 4471
rect 31726 4468 31754 4508
rect 32401 4505 32413 4508
rect 32447 4505 32459 4539
rect 32401 4499 32459 4505
rect 31527 4440 31754 4468
rect 31527 4437 31539 4440
rect 31481 4431 31539 4437
rect 31846 4428 31852 4480
rect 31904 4468 31910 4480
rect 32508 4468 32536 4635
rect 32582 4632 32588 4684
rect 32640 4672 32646 4684
rect 32640 4644 37872 4672
rect 32640 4632 32646 4644
rect 32677 4607 32735 4613
rect 32677 4573 32689 4607
rect 32723 4573 32735 4607
rect 32677 4567 32735 4573
rect 32692 4536 32720 4567
rect 33502 4564 33508 4616
rect 33560 4604 33566 4616
rect 33781 4607 33839 4613
rect 33781 4604 33793 4607
rect 33560 4576 33793 4604
rect 33560 4564 33566 4576
rect 33781 4573 33793 4576
rect 33827 4573 33839 4607
rect 33781 4567 33839 4573
rect 34330 4564 34336 4616
rect 34388 4604 34394 4616
rect 34698 4604 34704 4616
rect 34388 4576 34560 4604
rect 34659 4576 34704 4604
rect 34388 4564 34394 4576
rect 34422 4536 34428 4548
rect 32692 4508 34428 4536
rect 34422 4496 34428 4508
rect 34480 4496 34486 4548
rect 34532 4536 34560 4576
rect 34698 4564 34704 4576
rect 34756 4564 34762 4616
rect 35066 4604 35072 4616
rect 35027 4576 35072 4604
rect 35066 4564 35072 4576
rect 35124 4564 35130 4616
rect 35250 4564 35256 4616
rect 35308 4604 35314 4616
rect 37844 4613 37872 4644
rect 35897 4607 35955 4613
rect 35897 4604 35909 4607
rect 35308 4576 35909 4604
rect 35308 4564 35314 4576
rect 35897 4573 35909 4576
rect 35943 4573 35955 4607
rect 35897 4567 35955 4573
rect 37369 4607 37427 4613
rect 37369 4573 37381 4607
rect 37415 4573 37427 4607
rect 37369 4567 37427 4573
rect 37829 4607 37887 4613
rect 37829 4573 37841 4607
rect 37875 4573 37887 4607
rect 37829 4567 37887 4573
rect 34885 4539 34943 4545
rect 34885 4536 34897 4539
rect 34532 4508 34897 4536
rect 34885 4505 34897 4508
rect 34931 4505 34943 4539
rect 34885 4499 34943 4505
rect 34977 4539 35035 4545
rect 34977 4505 34989 4539
rect 35023 4536 35035 4539
rect 36538 4536 36544 4548
rect 35023 4508 36544 4536
rect 35023 4505 35035 4508
rect 34977 4499 35035 4505
rect 36538 4496 36544 4508
rect 36596 4496 36602 4548
rect 37384 4536 37412 4567
rect 37918 4536 37924 4548
rect 37384 4508 37924 4536
rect 37918 4496 37924 4508
rect 37976 4496 37982 4548
rect 31904 4440 32536 4468
rect 31904 4428 31910 4440
rect 34514 4428 34520 4480
rect 34572 4468 34578 4480
rect 35253 4471 35311 4477
rect 35253 4468 35265 4471
rect 34572 4440 35265 4468
rect 34572 4428 34578 4440
rect 35253 4437 35265 4440
rect 35299 4437 35311 4471
rect 35253 4431 35311 4437
rect 38013 4471 38071 4477
rect 38013 4437 38025 4471
rect 38059 4468 38071 4471
rect 38654 4468 38660 4480
rect 38059 4440 38660 4468
rect 38059 4437 38071 4440
rect 38013 4431 38071 4437
rect 38654 4428 38660 4440
rect 38712 4428 38718 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 11977 4267 12035 4273
rect 11977 4233 11989 4267
rect 12023 4264 12035 4267
rect 15194 4264 15200 4276
rect 12023 4236 15200 4264
rect 12023 4233 12035 4236
rect 11977 4227 12035 4233
rect 15194 4224 15200 4236
rect 15252 4224 15258 4276
rect 15286 4224 15292 4276
rect 15344 4264 15350 4276
rect 17770 4264 17776 4276
rect 15344 4236 17776 4264
rect 15344 4224 15350 4236
rect 8840 4199 8898 4205
rect 8840 4165 8852 4199
rect 8886 4196 8898 4199
rect 9122 4196 9128 4208
rect 8886 4168 9128 4196
rect 8886 4165 8898 4168
rect 8840 4159 8898 4165
rect 9122 4156 9128 4168
rect 9180 4156 9186 4208
rect 11514 4196 11520 4208
rect 11475 4168 11520 4196
rect 11514 4156 11520 4168
rect 11572 4156 11578 4208
rect 12802 4196 12808 4208
rect 12763 4168 12808 4196
rect 12802 4156 12808 4168
rect 12860 4156 12866 4208
rect 14274 4156 14280 4208
rect 14332 4196 14338 4208
rect 15381 4199 15439 4205
rect 15381 4196 15393 4199
rect 14332 4168 15393 4196
rect 14332 4156 14338 4168
rect 15381 4165 15393 4168
rect 15427 4165 15439 4199
rect 16298 4196 16304 4208
rect 15381 4159 15439 4165
rect 15488 4168 16304 4196
rect 8478 4088 8484 4140
rect 8536 4128 8542 4140
rect 8573 4131 8631 4137
rect 8573 4128 8585 4131
rect 8536 4100 8585 4128
rect 8536 4088 8542 4100
rect 8573 4097 8585 4100
rect 8619 4097 8631 4131
rect 8573 4091 8631 4097
rect 9582 4088 9588 4140
rect 9640 4128 9646 4140
rect 10781 4131 10839 4137
rect 9640 4100 10732 4128
rect 9640 4088 9646 4100
rect 10704 4069 10732 4100
rect 10781 4097 10793 4131
rect 10827 4128 10839 4131
rect 11330 4128 11336 4140
rect 10827 4100 11336 4128
rect 10827 4097 10839 4100
rect 10781 4091 10839 4097
rect 11330 4088 11336 4100
rect 11388 4088 11394 4140
rect 11793 4131 11851 4137
rect 11793 4097 11805 4131
rect 11839 4128 11851 4131
rect 12526 4128 12532 4140
rect 11839 4100 12532 4128
rect 11839 4097 11851 4100
rect 11793 4091 11851 4097
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 12713 4131 12771 4137
rect 12713 4097 12725 4131
rect 12759 4097 12771 4131
rect 12713 4091 12771 4097
rect 12897 4131 12955 4137
rect 12897 4097 12909 4131
rect 12943 4128 12955 4131
rect 13906 4128 13912 4140
rect 12943 4100 13768 4128
rect 13867 4100 13912 4128
rect 12943 4097 12955 4100
rect 12897 4091 12955 4097
rect 10597 4063 10655 4069
rect 10597 4060 10609 4063
rect 9968 4032 10609 4060
rect 9968 4001 9996 4032
rect 10597 4029 10609 4032
rect 10643 4029 10655 4063
rect 10597 4023 10655 4029
rect 10689 4063 10747 4069
rect 10689 4029 10701 4063
rect 10735 4029 10747 4063
rect 10689 4023 10747 4029
rect 9953 3995 10011 4001
rect 9953 3961 9965 3995
rect 9999 3961 10011 3995
rect 10410 3992 10416 4004
rect 10371 3964 10416 3992
rect 9953 3955 10011 3961
rect 10410 3952 10416 3964
rect 10468 3952 10474 4004
rect 10612 3992 10640 4023
rect 11146 4020 11152 4072
rect 11204 4060 11210 4072
rect 11609 4063 11667 4069
rect 11609 4060 11621 4063
rect 11204 4032 11621 4060
rect 11204 4020 11210 4032
rect 11609 4029 11621 4032
rect 11655 4029 11667 4063
rect 11609 4023 11667 4029
rect 11698 4020 11704 4072
rect 11756 4060 11762 4072
rect 12728 4060 12756 4091
rect 13740 4060 13768 4100
rect 13906 4088 13912 4100
rect 13964 4088 13970 4140
rect 14093 4131 14151 4137
rect 14093 4097 14105 4131
rect 14139 4097 14151 4131
rect 14642 4128 14648 4140
rect 14603 4100 14648 4128
rect 14093 4091 14151 4097
rect 13814 4060 13820 4072
rect 11756 4032 13216 4060
rect 13740 4032 13820 4060
rect 11756 4020 11762 4032
rect 10612 3964 11560 3992
rect 1670 3884 1676 3936
rect 1728 3924 1734 3936
rect 1949 3927 2007 3933
rect 1949 3924 1961 3927
rect 1728 3896 1961 3924
rect 1728 3884 1734 3896
rect 1949 3893 1961 3896
rect 1995 3893 2007 3927
rect 1949 3887 2007 3893
rect 3050 3884 3056 3936
rect 3108 3924 3114 3936
rect 8846 3924 8852 3936
rect 3108 3896 8852 3924
rect 3108 3884 3114 3896
rect 8846 3884 8852 3896
rect 8904 3884 8910 3936
rect 8938 3884 8944 3936
rect 8996 3924 9002 3936
rect 10428 3924 10456 3952
rect 10594 3924 10600 3936
rect 8996 3896 10456 3924
rect 10555 3896 10600 3924
rect 8996 3884 9002 3896
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 11532 3933 11560 3964
rect 11517 3927 11575 3933
rect 11517 3893 11529 3927
rect 11563 3893 11575 3927
rect 11517 3887 11575 3893
rect 12710 3884 12716 3936
rect 12768 3924 12774 3936
rect 13081 3927 13139 3933
rect 13081 3924 13093 3927
rect 12768 3896 13093 3924
rect 12768 3884 12774 3896
rect 13081 3893 13093 3896
rect 13127 3893 13139 3927
rect 13188 3924 13216 4032
rect 13814 4020 13820 4032
rect 13872 4020 13878 4072
rect 13998 4060 14004 4072
rect 13959 4032 14004 4060
rect 13998 4020 14004 4032
rect 14056 4020 14062 4072
rect 14108 4060 14136 4091
rect 14642 4088 14648 4100
rect 14700 4088 14706 4140
rect 15488 4128 15516 4168
rect 16298 4156 16304 4168
rect 16356 4156 16362 4208
rect 15654 4128 15660 4140
rect 14844 4100 15516 4128
rect 15615 4100 15660 4128
rect 14844 4060 14872 4100
rect 15654 4088 15660 4100
rect 15712 4088 15718 4140
rect 16853 4131 16911 4137
rect 16853 4097 16865 4131
rect 16899 4128 16911 4131
rect 17034 4128 17040 4140
rect 16899 4100 17040 4128
rect 16899 4097 16911 4100
rect 16853 4091 16911 4097
rect 17034 4088 17040 4100
rect 17092 4088 17098 4140
rect 17236 4128 17264 4236
rect 17770 4224 17776 4236
rect 17828 4224 17834 4276
rect 19150 4224 19156 4276
rect 19208 4264 19214 4276
rect 19429 4267 19487 4273
rect 19429 4264 19441 4267
rect 19208 4236 19441 4264
rect 19208 4224 19214 4236
rect 19429 4233 19441 4236
rect 19475 4233 19487 4267
rect 21082 4264 21088 4276
rect 19429 4227 19487 4233
rect 20272 4236 21088 4264
rect 18230 4156 18236 4208
rect 18288 4196 18294 4208
rect 20272 4205 20300 4236
rect 21082 4224 21088 4236
rect 21140 4224 21146 4276
rect 22002 4224 22008 4276
rect 22060 4264 22066 4276
rect 23201 4267 23259 4273
rect 23201 4264 23213 4267
rect 22060 4236 23213 4264
rect 22060 4224 22066 4236
rect 23201 4233 23213 4236
rect 23247 4264 23259 4267
rect 24394 4264 24400 4276
rect 23247 4236 24400 4264
rect 23247 4233 23259 4236
rect 23201 4227 23259 4233
rect 24394 4224 24400 4236
rect 24452 4224 24458 4276
rect 29546 4224 29552 4276
rect 29604 4264 29610 4276
rect 31202 4264 31208 4276
rect 29604 4236 31208 4264
rect 29604 4224 29610 4236
rect 18969 4199 19027 4205
rect 18969 4196 18981 4199
rect 18288 4168 18981 4196
rect 18288 4156 18294 4168
rect 18969 4165 18981 4168
rect 19015 4165 19027 4199
rect 20257 4199 20315 4205
rect 18969 4159 19027 4165
rect 19076 4168 19380 4196
rect 17313 4131 17371 4137
rect 17313 4128 17325 4131
rect 17236 4100 17325 4128
rect 17313 4097 17325 4100
rect 17359 4097 17371 4131
rect 17313 4091 17371 4097
rect 17681 4131 17739 4137
rect 17681 4097 17693 4131
rect 17727 4128 17739 4131
rect 18046 4128 18052 4140
rect 17727 4100 18052 4128
rect 17727 4097 17739 4100
rect 17681 4091 17739 4097
rect 18046 4088 18052 4100
rect 18104 4088 18110 4140
rect 18325 4131 18383 4137
rect 18325 4097 18337 4131
rect 18371 4097 18383 4131
rect 18325 4091 18383 4097
rect 14108 4032 14872 4060
rect 14918 4020 14924 4072
rect 14976 4060 14982 4072
rect 15473 4063 15531 4069
rect 15473 4060 15485 4063
rect 14976 4032 15485 4060
rect 14976 4020 14982 4032
rect 15473 4029 15485 4032
rect 15519 4029 15531 4063
rect 16758 4060 16764 4072
rect 15473 4023 15531 4029
rect 15580 4032 16764 4060
rect 13630 3952 13636 4004
rect 13688 3992 13694 4004
rect 15580 3992 15608 4032
rect 16758 4020 16764 4032
rect 16816 4020 16822 4072
rect 17497 4063 17555 4069
rect 17497 4029 17509 4063
rect 17543 4060 17555 4063
rect 18230 4060 18236 4072
rect 17543 4032 18236 4060
rect 17543 4029 17555 4032
rect 17497 4023 17555 4029
rect 18230 4020 18236 4032
rect 18288 4020 18294 4072
rect 13688 3964 15608 3992
rect 15841 3995 15899 4001
rect 13688 3952 13694 3964
rect 15841 3961 15853 3995
rect 15887 3992 15899 3995
rect 16390 3992 16396 4004
rect 15887 3964 16396 3992
rect 15887 3961 15899 3964
rect 15841 3955 15899 3961
rect 16390 3952 16396 3964
rect 16448 3952 16454 4004
rect 17586 3992 17592 4004
rect 17547 3964 17592 3992
rect 17586 3952 17592 3964
rect 17644 3952 17650 4004
rect 17770 3952 17776 4004
rect 17828 3992 17834 4004
rect 18340 3992 18368 4091
rect 18506 4088 18512 4140
rect 18564 4128 18570 4140
rect 19076 4128 19104 4168
rect 19242 4128 19248 4140
rect 18564 4100 19104 4128
rect 19203 4100 19248 4128
rect 18564 4088 18570 4100
rect 19242 4088 19248 4100
rect 19300 4088 19306 4140
rect 19352 4128 19380 4168
rect 20257 4165 20269 4199
rect 20303 4165 20315 4199
rect 20257 4159 20315 4165
rect 22088 4199 22146 4205
rect 22088 4165 22100 4199
rect 22134 4196 22146 4199
rect 22186 4196 22192 4208
rect 22134 4168 22192 4196
rect 22134 4165 22146 4168
rect 22088 4159 22146 4165
rect 22186 4156 22192 4168
rect 22244 4156 22250 4208
rect 24029 4199 24087 4205
rect 24029 4165 24041 4199
rect 24075 4196 24087 4199
rect 24762 4196 24768 4208
rect 24075 4168 24768 4196
rect 24075 4165 24087 4168
rect 24029 4159 24087 4165
rect 24762 4156 24768 4168
rect 24820 4156 24826 4208
rect 26234 4156 26240 4208
rect 26292 4196 26298 4208
rect 29365 4199 29423 4205
rect 29365 4196 29377 4199
rect 26292 4168 29377 4196
rect 26292 4156 26298 4168
rect 29365 4165 29377 4168
rect 29411 4165 29423 4199
rect 30374 4196 30380 4208
rect 29365 4159 29423 4165
rect 29564 4168 30380 4196
rect 21082 4128 21088 4140
rect 19352 4100 20484 4128
rect 21043 4100 21088 4128
rect 19150 4060 19156 4072
rect 19111 4032 19156 4060
rect 19150 4020 19156 4032
rect 19208 4020 19214 4072
rect 20346 4060 20352 4072
rect 19260 4032 20352 4060
rect 17828 3964 18368 3992
rect 17828 3952 17834 3964
rect 14458 3924 14464 3936
rect 13188 3896 14464 3924
rect 13081 3887 13139 3893
rect 14458 3884 14464 3896
rect 14516 3884 14522 3936
rect 14829 3927 14887 3933
rect 14829 3893 14841 3927
rect 14875 3924 14887 3927
rect 15286 3924 15292 3936
rect 14875 3896 15292 3924
rect 14875 3893 14887 3896
rect 14829 3887 14887 3893
rect 15286 3884 15292 3896
rect 15344 3884 15350 3936
rect 15470 3924 15476 3936
rect 15431 3896 15476 3924
rect 15470 3884 15476 3896
rect 15528 3884 15534 3936
rect 16666 3924 16672 3936
rect 16627 3896 16672 3924
rect 16666 3884 16672 3896
rect 16724 3884 16730 3936
rect 17218 3884 17224 3936
rect 17276 3924 17282 3936
rect 17497 3927 17555 3933
rect 17497 3924 17509 3927
rect 17276 3896 17509 3924
rect 17276 3884 17282 3896
rect 17497 3893 17509 3896
rect 17543 3893 17555 3927
rect 17497 3887 17555 3893
rect 17678 3884 17684 3936
rect 17736 3924 17742 3936
rect 19260 3933 19288 4032
rect 20346 4020 20352 4032
rect 20404 4020 20410 4072
rect 20456 4060 20484 4100
rect 21082 4088 21088 4100
rect 21140 4088 21146 4140
rect 24486 4088 24492 4140
rect 24544 4128 24550 4140
rect 24949 4131 25007 4137
rect 24949 4128 24961 4131
rect 24544 4100 24961 4128
rect 24544 4088 24550 4100
rect 24949 4097 24961 4100
rect 24995 4097 25007 4131
rect 25958 4128 25964 4140
rect 25919 4100 25964 4128
rect 24949 4091 25007 4097
rect 25958 4088 25964 4100
rect 26016 4088 26022 4140
rect 26973 4131 27031 4137
rect 26973 4097 26985 4131
rect 27019 4128 27031 4131
rect 27154 4128 27160 4140
rect 27019 4100 27160 4128
rect 27019 4097 27031 4100
rect 26973 4091 27031 4097
rect 27154 4088 27160 4100
rect 27212 4088 27218 4140
rect 27338 4088 27344 4140
rect 27396 4128 27402 4140
rect 27709 4131 27767 4137
rect 27709 4128 27721 4131
rect 27396 4100 27721 4128
rect 27396 4088 27402 4100
rect 27709 4097 27721 4100
rect 27755 4097 27767 4131
rect 27709 4091 27767 4097
rect 28629 4131 28687 4137
rect 28629 4097 28641 4131
rect 28675 4097 28687 4131
rect 29564 4128 29592 4168
rect 30374 4156 30380 4168
rect 30432 4156 30438 4208
rect 30576 4205 30604 4236
rect 31202 4224 31208 4236
rect 31260 4224 31266 4276
rect 32030 4224 32036 4276
rect 32088 4264 32094 4276
rect 34330 4264 34336 4276
rect 32088 4236 34336 4264
rect 32088 4224 32094 4236
rect 34330 4224 34336 4236
rect 34388 4224 34394 4276
rect 34606 4224 34612 4276
rect 34664 4264 34670 4276
rect 34701 4267 34759 4273
rect 34701 4264 34713 4267
rect 34664 4236 34713 4264
rect 34664 4224 34670 4236
rect 34701 4233 34713 4236
rect 34747 4233 34759 4267
rect 34701 4227 34759 4233
rect 35066 4224 35072 4276
rect 35124 4264 35130 4276
rect 35434 4264 35440 4276
rect 35124 4236 35440 4264
rect 35124 4224 35130 4236
rect 35434 4224 35440 4236
rect 35492 4224 35498 4276
rect 36538 4264 36544 4276
rect 36499 4236 36544 4264
rect 36538 4224 36544 4236
rect 36596 4224 36602 4276
rect 30561 4199 30619 4205
rect 30561 4165 30573 4199
rect 30607 4165 30619 4199
rect 31110 4196 31116 4208
rect 30561 4159 30619 4165
rect 30852 4168 31116 4196
rect 28629 4091 28687 4097
rect 28736 4100 29592 4128
rect 29641 4131 29699 4137
rect 21450 4060 21456 4072
rect 20456 4032 21456 4060
rect 21450 4020 21456 4032
rect 21508 4020 21514 4072
rect 21821 4063 21879 4069
rect 21821 4029 21833 4063
rect 21867 4029 21879 4063
rect 21821 4023 21879 4029
rect 24673 4063 24731 4069
rect 24673 4029 24685 4063
rect 24719 4060 24731 4063
rect 24719 4032 24992 4060
rect 24719 4029 24731 4032
rect 24673 4023 24731 4029
rect 19610 3952 19616 4004
rect 19668 3992 19674 4004
rect 20070 3992 20076 4004
rect 19668 3964 20076 3992
rect 19668 3952 19674 3964
rect 20070 3952 20076 3964
rect 20128 3952 20134 4004
rect 21726 3992 21732 4004
rect 20180 3964 21732 3992
rect 18141 3927 18199 3933
rect 18141 3924 18153 3927
rect 17736 3896 18153 3924
rect 17736 3884 17742 3896
rect 18141 3893 18153 3896
rect 18187 3893 18199 3927
rect 18141 3887 18199 3893
rect 19245 3927 19303 3933
rect 19245 3893 19257 3927
rect 19291 3893 19303 3927
rect 19245 3887 19303 3893
rect 19518 3884 19524 3936
rect 19576 3924 19582 3936
rect 20180 3924 20208 3964
rect 21726 3952 21732 3964
rect 21784 3952 21790 4004
rect 20346 3924 20352 3936
rect 19576 3896 20208 3924
rect 20307 3896 20352 3924
rect 19576 3884 19582 3896
rect 20346 3884 20352 3896
rect 20404 3884 20410 3936
rect 20898 3924 20904 3936
rect 20859 3896 20904 3924
rect 20898 3884 20904 3896
rect 20956 3884 20962 3936
rect 21836 3924 21864 4023
rect 24964 4004 24992 4032
rect 25682 4020 25688 4072
rect 25740 4060 25746 4072
rect 28644 4060 28672 4091
rect 25740 4032 28672 4060
rect 25740 4020 25746 4032
rect 24213 3995 24271 4001
rect 24213 3961 24225 3995
rect 24259 3992 24271 3995
rect 24854 3992 24860 4004
rect 24259 3964 24860 3992
rect 24259 3961 24271 3964
rect 24213 3955 24271 3961
rect 24854 3952 24860 3964
rect 24912 3952 24918 4004
rect 24946 3952 24952 4004
rect 25004 3952 25010 4004
rect 25332 3964 27292 3992
rect 22094 3924 22100 3936
rect 21836 3896 22100 3924
rect 22094 3884 22100 3896
rect 22152 3884 22158 3936
rect 22554 3884 22560 3936
rect 22612 3924 22618 3936
rect 25332 3924 25360 3964
rect 22612 3896 25360 3924
rect 22612 3884 22618 3896
rect 25406 3884 25412 3936
rect 25464 3924 25470 3936
rect 26145 3927 26203 3933
rect 26145 3924 26157 3927
rect 25464 3896 26157 3924
rect 25464 3884 25470 3896
rect 26145 3893 26157 3896
rect 26191 3893 26203 3927
rect 26145 3887 26203 3893
rect 26418 3884 26424 3936
rect 26476 3924 26482 3936
rect 27157 3927 27215 3933
rect 27157 3924 27169 3927
rect 26476 3896 27169 3924
rect 26476 3884 26482 3896
rect 27157 3893 27169 3896
rect 27203 3893 27215 3927
rect 27264 3924 27292 3964
rect 27338 3952 27344 4004
rect 27396 3992 27402 4004
rect 28445 3995 28503 4001
rect 28445 3992 28457 3995
rect 27396 3964 28457 3992
rect 27396 3952 27402 3964
rect 28445 3961 28457 3964
rect 28491 3961 28503 3995
rect 28445 3955 28503 3961
rect 27522 3924 27528 3936
rect 27264 3896 27528 3924
rect 27157 3887 27215 3893
rect 27522 3884 27528 3896
rect 27580 3884 27586 3936
rect 27614 3884 27620 3936
rect 27672 3924 27678 3936
rect 27893 3927 27951 3933
rect 27893 3924 27905 3927
rect 27672 3896 27905 3924
rect 27672 3884 27678 3896
rect 27893 3893 27905 3896
rect 27939 3893 27951 3927
rect 27893 3887 27951 3893
rect 28350 3884 28356 3936
rect 28408 3924 28414 3936
rect 28736 3924 28764 4100
rect 29641 4097 29653 4131
rect 29687 4128 29699 4131
rect 30852 4128 30880 4168
rect 31110 4156 31116 4168
rect 31168 4156 31174 4208
rect 31662 4156 31668 4208
rect 31720 4196 31726 4208
rect 36170 4196 36176 4208
rect 31720 4168 36176 4196
rect 31720 4156 31726 4168
rect 36170 4156 36176 4168
rect 36228 4156 36234 4208
rect 29687 4100 30880 4128
rect 30929 4131 30987 4137
rect 29687 4097 29699 4100
rect 29641 4091 29699 4097
rect 30929 4097 30941 4131
rect 30975 4128 30987 4131
rect 30975 4100 31340 4128
rect 30975 4097 30987 4100
rect 30929 4091 30987 4097
rect 29454 4060 29460 4072
rect 29415 4032 29460 4060
rect 29454 4020 29460 4032
rect 29512 4020 29518 4072
rect 29546 4020 29552 4072
rect 29604 4060 29610 4072
rect 30742 4060 30748 4072
rect 29604 4032 30512 4060
rect 30703 4032 30748 4060
rect 29604 4020 29610 4032
rect 30374 3992 30380 4004
rect 29656 3964 30380 3992
rect 29656 3933 29684 3964
rect 30374 3952 30380 3964
rect 30432 3952 30438 4004
rect 30484 3992 30512 4032
rect 30742 4020 30748 4032
rect 30800 4020 30806 4072
rect 30837 4063 30895 4069
rect 30837 4029 30849 4063
rect 30883 4060 30895 4063
rect 31202 4060 31208 4072
rect 30883 4032 31208 4060
rect 30883 4029 30895 4032
rect 30837 4023 30895 4029
rect 31202 4020 31208 4032
rect 31260 4020 31266 4072
rect 31312 3992 31340 4100
rect 31386 4088 31392 4140
rect 31444 4128 31450 4140
rect 31573 4131 31631 4137
rect 31573 4128 31585 4131
rect 31444 4100 31585 4128
rect 31444 4088 31450 4100
rect 31573 4097 31585 4100
rect 31619 4097 31631 4131
rect 32306 4128 32312 4140
rect 32267 4100 32312 4128
rect 31573 4091 31631 4097
rect 32306 4088 32312 4100
rect 32364 4088 32370 4140
rect 32953 4131 33011 4137
rect 32953 4097 32965 4131
rect 32999 4097 33011 4131
rect 32953 4091 33011 4097
rect 33597 4131 33655 4137
rect 33597 4097 33609 4131
rect 33643 4097 33655 4131
rect 34514 4128 34520 4140
rect 34475 4100 34520 4128
rect 33597 4091 33655 4097
rect 31662 4020 31668 4072
rect 31720 4060 31726 4072
rect 32968 4060 32996 4091
rect 31720 4032 32996 4060
rect 31720 4020 31726 4032
rect 32769 3995 32827 4001
rect 32769 3992 32781 3995
rect 30484 3964 30880 3992
rect 31312 3964 32781 3992
rect 28408 3896 28764 3924
rect 29641 3927 29699 3933
rect 28408 3884 28414 3896
rect 29641 3893 29653 3927
rect 29687 3893 29699 3927
rect 29822 3924 29828 3936
rect 29783 3896 29828 3924
rect 29641 3887 29699 3893
rect 29822 3884 29828 3896
rect 29880 3884 29886 3936
rect 30466 3884 30472 3936
rect 30524 3924 30530 3936
rect 30745 3927 30803 3933
rect 30745 3924 30757 3927
rect 30524 3896 30757 3924
rect 30524 3884 30530 3896
rect 30745 3893 30757 3896
rect 30791 3893 30803 3927
rect 30852 3924 30880 3964
rect 32769 3961 32781 3964
rect 32815 3961 32827 3995
rect 33612 3992 33640 4091
rect 34514 4088 34520 4100
rect 34572 4088 34578 4140
rect 34606 4088 34612 4140
rect 34664 4128 34670 4140
rect 35345 4131 35403 4137
rect 35345 4128 35357 4131
rect 34664 4100 35357 4128
rect 34664 4088 34670 4100
rect 35345 4097 35357 4100
rect 35391 4097 35403 4131
rect 35345 4091 35403 4097
rect 35802 4088 35808 4140
rect 35860 4128 35866 4140
rect 35989 4131 36047 4137
rect 35989 4128 36001 4131
rect 35860 4100 36001 4128
rect 35860 4088 35866 4100
rect 35989 4097 36001 4100
rect 36035 4097 36047 4131
rect 35989 4091 36047 4097
rect 36725 4131 36783 4137
rect 36725 4097 36737 4131
rect 36771 4128 36783 4131
rect 36814 4128 36820 4140
rect 36771 4100 36820 4128
rect 36771 4097 36783 4100
rect 36725 4091 36783 4097
rect 36814 4088 36820 4100
rect 36872 4088 36878 4140
rect 37642 4128 37648 4140
rect 37603 4100 37648 4128
rect 37642 4088 37648 4100
rect 37700 4088 37706 4140
rect 33778 4020 33784 4072
rect 33836 4060 33842 4072
rect 34333 4063 34391 4069
rect 34333 4060 34345 4063
rect 33836 4032 34345 4060
rect 33836 4020 33842 4032
rect 34333 4029 34345 4032
rect 34379 4029 34391 4063
rect 34333 4023 34391 4029
rect 32769 3955 32827 3961
rect 32876 3964 33640 3992
rect 31389 3927 31447 3933
rect 31389 3924 31401 3927
rect 30852 3896 31401 3924
rect 30745 3887 30803 3893
rect 31389 3893 31401 3896
rect 31435 3893 31447 3927
rect 31389 3887 31447 3893
rect 31478 3884 31484 3936
rect 31536 3924 31542 3936
rect 32125 3927 32183 3933
rect 32125 3924 32137 3927
rect 31536 3896 32137 3924
rect 31536 3884 31542 3896
rect 32125 3893 32137 3896
rect 32171 3893 32183 3927
rect 32125 3887 32183 3893
rect 32398 3884 32404 3936
rect 32456 3924 32462 3936
rect 32876 3924 32904 3964
rect 33870 3952 33876 4004
rect 33928 3992 33934 4004
rect 35250 3992 35256 4004
rect 33928 3964 35256 3992
rect 33928 3952 33934 3964
rect 35250 3952 35256 3964
rect 35308 3952 35314 4004
rect 35618 3952 35624 4004
rect 35676 3992 35682 4004
rect 35805 3995 35863 4001
rect 35805 3992 35817 3995
rect 35676 3964 35817 3992
rect 35676 3952 35682 3964
rect 35805 3961 35817 3964
rect 35851 3961 35863 3995
rect 35805 3955 35863 3961
rect 32456 3896 32904 3924
rect 32456 3884 32462 3896
rect 32950 3884 32956 3936
rect 33008 3924 33014 3936
rect 33413 3927 33471 3933
rect 33413 3924 33425 3927
rect 33008 3896 33425 3924
rect 33008 3884 33014 3896
rect 33413 3893 33425 3896
rect 33459 3893 33471 3927
rect 33413 3887 33471 3893
rect 34790 3884 34796 3936
rect 34848 3924 34854 3936
rect 35161 3927 35219 3933
rect 35161 3924 35173 3927
rect 34848 3896 35173 3924
rect 34848 3884 34854 3896
rect 35161 3893 35173 3896
rect 35207 3893 35219 3927
rect 35161 3887 35219 3893
rect 37550 3884 37556 3936
rect 37608 3924 37614 3936
rect 37829 3927 37887 3933
rect 37829 3924 37841 3927
rect 37608 3896 37841 3924
rect 37608 3884 37614 3896
rect 37829 3893 37841 3896
rect 37875 3893 37887 3927
rect 37829 3887 37887 3893
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 3789 3723 3847 3729
rect 3789 3689 3801 3723
rect 3835 3720 3847 3723
rect 4614 3720 4620 3732
rect 3835 3692 4620 3720
rect 3835 3689 3847 3692
rect 3789 3683 3847 3689
rect 4614 3680 4620 3692
rect 4672 3680 4678 3732
rect 6549 3723 6607 3729
rect 6549 3689 6561 3723
rect 6595 3720 6607 3723
rect 8110 3720 8116 3732
rect 6595 3692 8116 3720
rect 6595 3689 6607 3692
rect 6549 3683 6607 3689
rect 8110 3680 8116 3692
rect 8168 3680 8174 3732
rect 9125 3723 9183 3729
rect 9125 3720 9137 3723
rect 8220 3692 9137 3720
rect 7558 3652 7564 3664
rect 7519 3624 7564 3652
rect 7558 3612 7564 3624
rect 7616 3612 7622 3664
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 1581 3519 1639 3525
rect 1581 3516 1593 3519
rect 1360 3488 1593 3516
rect 1360 3476 1366 3488
rect 1581 3485 1593 3488
rect 1627 3485 1639 3519
rect 1581 3479 1639 3485
rect 2406 3476 2412 3528
rect 2464 3516 2470 3528
rect 2685 3519 2743 3525
rect 2685 3516 2697 3519
rect 2464 3488 2697 3516
rect 2464 3476 2470 3488
rect 2685 3485 2697 3488
rect 2731 3485 2743 3519
rect 2685 3479 2743 3485
rect 3510 3476 3516 3528
rect 3568 3516 3574 3528
rect 3973 3519 4031 3525
rect 3973 3516 3985 3519
rect 3568 3488 3985 3516
rect 3568 3476 3574 3488
rect 3973 3485 3985 3488
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 6733 3519 6791 3525
rect 6733 3516 6745 3519
rect 6512 3488 6745 3516
rect 6512 3476 6518 3488
rect 6733 3485 6745 3488
rect 6779 3485 6791 3519
rect 6733 3479 6791 3485
rect 7745 3519 7803 3525
rect 7745 3485 7757 3519
rect 7791 3516 7803 3519
rect 7926 3516 7932 3528
rect 7791 3488 7932 3516
rect 7791 3485 7803 3488
rect 7745 3479 7803 3485
rect 7926 3476 7932 3488
rect 7984 3476 7990 3528
rect 8220 3525 8248 3692
rect 9125 3689 9137 3692
rect 9171 3689 9183 3723
rect 9125 3683 9183 3689
rect 9217 3723 9275 3729
rect 9217 3689 9229 3723
rect 9263 3720 9275 3723
rect 9582 3720 9588 3732
rect 9263 3692 9588 3720
rect 9263 3689 9275 3692
rect 9217 3683 9275 3689
rect 9582 3680 9588 3692
rect 9640 3680 9646 3732
rect 11146 3720 11152 3732
rect 11107 3692 11152 3720
rect 11146 3680 11152 3692
rect 11204 3680 11210 3732
rect 12526 3680 12532 3732
rect 12584 3720 12590 3732
rect 12989 3723 13047 3729
rect 12989 3720 13001 3723
rect 12584 3692 13001 3720
rect 12584 3680 12590 3692
rect 12989 3689 13001 3692
rect 13035 3689 13047 3723
rect 12989 3683 13047 3689
rect 14182 3680 14188 3732
rect 14240 3720 14246 3732
rect 14461 3723 14519 3729
rect 14461 3720 14473 3723
rect 14240 3692 14473 3720
rect 14240 3680 14246 3692
rect 14461 3689 14473 3692
rect 14507 3689 14519 3723
rect 14461 3683 14519 3689
rect 15654 3680 15660 3732
rect 15712 3720 15718 3732
rect 16758 3720 16764 3732
rect 15712 3692 16764 3720
rect 15712 3680 15718 3692
rect 16758 3680 16764 3692
rect 16816 3720 16822 3732
rect 16853 3723 16911 3729
rect 16853 3720 16865 3723
rect 16816 3692 16865 3720
rect 16816 3680 16822 3692
rect 16853 3689 16865 3692
rect 16899 3689 16911 3723
rect 16853 3683 16911 3689
rect 16942 3680 16948 3732
rect 17000 3720 17006 3732
rect 17313 3723 17371 3729
rect 17313 3720 17325 3723
rect 17000 3692 17325 3720
rect 17000 3680 17006 3692
rect 17313 3689 17325 3692
rect 17359 3689 17371 3723
rect 17313 3683 17371 3689
rect 19242 3680 19248 3732
rect 19300 3720 19306 3732
rect 20714 3720 20720 3732
rect 19300 3692 20720 3720
rect 19300 3680 19306 3692
rect 20714 3680 20720 3692
rect 20772 3720 20778 3732
rect 21361 3723 21419 3729
rect 21361 3720 21373 3723
rect 20772 3692 21373 3720
rect 20772 3680 20778 3692
rect 21361 3689 21373 3692
rect 21407 3689 21419 3723
rect 21361 3683 21419 3689
rect 21450 3680 21456 3732
rect 21508 3720 21514 3732
rect 24578 3720 24584 3732
rect 21508 3692 24440 3720
rect 24539 3692 24584 3720
rect 21508 3680 21514 3692
rect 8478 3612 8484 3664
rect 8536 3652 8542 3664
rect 8536 3624 9812 3652
rect 8536 3612 8542 3624
rect 8938 3584 8944 3596
rect 8899 3556 8944 3584
rect 8938 3544 8944 3556
rect 8996 3544 9002 3596
rect 9122 3544 9128 3596
rect 9180 3584 9186 3596
rect 9628 3584 9634 3596
rect 9180 3556 9634 3584
rect 9180 3544 9186 3556
rect 9628 3544 9634 3556
rect 9686 3544 9692 3596
rect 9784 3593 9812 3624
rect 17126 3612 17132 3664
rect 17184 3652 17190 3664
rect 19886 3652 19892 3664
rect 17184 3624 19892 3652
rect 17184 3612 17190 3624
rect 19886 3612 19892 3624
rect 19944 3612 19950 3664
rect 23845 3655 23903 3661
rect 23845 3621 23857 3655
rect 23891 3621 23903 3655
rect 24412 3652 24440 3692
rect 24578 3680 24584 3692
rect 24636 3680 24642 3732
rect 24949 3723 25007 3729
rect 24949 3689 24961 3723
rect 24995 3720 25007 3723
rect 26234 3720 26240 3732
rect 24995 3692 26240 3720
rect 24995 3689 25007 3692
rect 24949 3683 25007 3689
rect 26234 3680 26240 3692
rect 26292 3680 26298 3732
rect 27154 3720 27160 3732
rect 27115 3692 27160 3720
rect 27154 3680 27160 3692
rect 27212 3680 27218 3732
rect 27246 3680 27252 3732
rect 27304 3720 27310 3732
rect 29914 3720 29920 3732
rect 27304 3692 29920 3720
rect 27304 3680 27310 3692
rect 29914 3680 29920 3692
rect 29972 3680 29978 3732
rect 30282 3680 30288 3732
rect 30340 3720 30346 3732
rect 32306 3720 32312 3732
rect 30340 3692 32312 3720
rect 30340 3680 30346 3692
rect 32306 3680 32312 3692
rect 32364 3680 32370 3732
rect 32766 3680 32772 3732
rect 32824 3720 32830 3732
rect 34054 3720 34060 3732
rect 32824 3692 34060 3720
rect 32824 3680 32830 3692
rect 34054 3680 34060 3692
rect 34112 3680 34118 3732
rect 29822 3652 29828 3664
rect 24412 3624 29828 3652
rect 23845 3615 23903 3621
rect 9758 3587 9816 3593
rect 9758 3553 9770 3587
rect 9804 3553 9816 3587
rect 9758 3547 9816 3553
rect 12986 3544 12992 3596
rect 13044 3584 13050 3596
rect 14093 3587 14151 3593
rect 14093 3584 14105 3587
rect 13044 3556 14105 3584
rect 13044 3544 13050 3556
rect 14093 3553 14105 3556
rect 14139 3553 14151 3587
rect 14093 3547 14151 3553
rect 16942 3544 16948 3596
rect 17000 3584 17006 3596
rect 17770 3584 17776 3596
rect 17000 3556 17776 3584
rect 17000 3544 17006 3556
rect 17770 3544 17776 3556
rect 17828 3544 17834 3596
rect 19058 3544 19064 3596
rect 19116 3584 19122 3596
rect 19610 3584 19616 3596
rect 19116 3556 19616 3584
rect 19116 3544 19122 3556
rect 19610 3544 19616 3556
rect 19668 3544 19674 3596
rect 22094 3584 22100 3596
rect 21284 3556 22100 3584
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3516 8447 3519
rect 9030 3516 9036 3528
rect 8435 3488 9036 3516
rect 8435 3485 8447 3488
rect 8389 3479 8447 3485
rect 9030 3476 9036 3488
rect 9088 3476 9094 3528
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3516 9367 3519
rect 9858 3516 9864 3528
rect 9355 3488 9864 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 9858 3476 9864 3488
rect 9916 3476 9922 3528
rect 10036 3519 10094 3525
rect 10036 3510 10048 3519
rect 9968 3485 10048 3510
rect 10082 3485 10094 3519
rect 9968 3482 10094 3485
rect 4614 3408 4620 3460
rect 4672 3448 4678 3460
rect 9766 3448 9772 3460
rect 4672 3420 9772 3448
rect 4672 3408 4678 3420
rect 9766 3408 9772 3420
rect 9824 3408 9830 3460
rect 9968 3448 9996 3482
rect 10036 3479 10094 3482
rect 11609 3519 11667 3525
rect 11609 3485 11621 3519
rect 11655 3516 11667 3519
rect 13538 3516 13544 3528
rect 11655 3488 13544 3516
rect 11655 3485 11667 3488
rect 11609 3479 11667 3485
rect 13538 3476 13544 3488
rect 13596 3476 13602 3528
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3516 14335 3519
rect 14826 3516 14832 3528
rect 14323 3488 14832 3516
rect 14323 3485 14335 3488
rect 14277 3479 14335 3485
rect 14826 3476 14832 3488
rect 14884 3476 14890 3528
rect 15473 3519 15531 3525
rect 15473 3485 15485 3519
rect 15519 3516 15531 3519
rect 16850 3516 16856 3528
rect 15519 3488 16856 3516
rect 15519 3485 15531 3488
rect 15473 3479 15531 3485
rect 16850 3476 16856 3488
rect 16908 3476 16914 3528
rect 17497 3519 17555 3525
rect 17497 3485 17509 3519
rect 17543 3485 17555 3519
rect 17497 3479 17555 3485
rect 18509 3519 18567 3525
rect 18509 3485 18521 3519
rect 18555 3516 18567 3519
rect 19426 3516 19432 3528
rect 18555 3488 19432 3516
rect 18555 3485 18567 3488
rect 18509 3479 18567 3485
rect 9876 3420 9996 3448
rect 11876 3451 11934 3457
rect 1397 3383 1455 3389
rect 1397 3349 1409 3383
rect 1443 3380 1455 3383
rect 2222 3380 2228 3392
rect 1443 3352 2228 3380
rect 1443 3349 1455 3352
rect 1397 3343 1455 3349
rect 2222 3340 2228 3352
rect 2280 3340 2286 3392
rect 2501 3383 2559 3389
rect 2501 3349 2513 3383
rect 2547 3380 2559 3383
rect 2866 3380 2872 3392
rect 2547 3352 2872 3380
rect 2547 3349 2559 3352
rect 2501 3343 2559 3349
rect 2866 3340 2872 3352
rect 2924 3340 2930 3392
rect 8294 3380 8300 3392
rect 8255 3352 8300 3380
rect 8294 3340 8300 3352
rect 8352 3340 8358 3392
rect 9674 3340 9680 3392
rect 9732 3380 9738 3392
rect 9876 3380 9904 3420
rect 11876 3417 11888 3451
rect 11922 3448 11934 3451
rect 12066 3448 12072 3460
rect 11922 3420 12072 3448
rect 11922 3417 11934 3420
rect 11876 3411 11934 3417
rect 12066 3408 12072 3420
rect 12124 3408 12130 3460
rect 15740 3451 15798 3457
rect 15740 3417 15752 3451
rect 15786 3448 15798 3451
rect 16666 3448 16672 3460
rect 15786 3420 16672 3448
rect 15786 3417 15798 3420
rect 15740 3411 15798 3417
rect 16666 3408 16672 3420
rect 16724 3408 16730 3460
rect 9732 3352 9904 3380
rect 9732 3340 9738 3352
rect 9950 3340 9956 3392
rect 10008 3380 10014 3392
rect 11054 3380 11060 3392
rect 10008 3352 11060 3380
rect 10008 3340 10014 3352
rect 11054 3340 11060 3352
rect 11112 3340 11118 3392
rect 13814 3340 13820 3392
rect 13872 3380 13878 3392
rect 14642 3380 14648 3392
rect 13872 3352 14648 3380
rect 13872 3340 13878 3352
rect 14642 3340 14648 3352
rect 14700 3340 14706 3392
rect 15838 3340 15844 3392
rect 15896 3380 15902 3392
rect 17512 3380 17540 3479
rect 19426 3476 19432 3488
rect 19484 3476 19490 3528
rect 19981 3519 20039 3525
rect 19981 3485 19993 3519
rect 20027 3516 20039 3519
rect 21284 3516 21312 3556
rect 22094 3544 22100 3556
rect 22152 3584 22158 3596
rect 22465 3587 22523 3593
rect 22465 3584 22477 3587
rect 22152 3556 22477 3584
rect 22152 3544 22158 3556
rect 22465 3553 22477 3556
rect 22511 3553 22523 3587
rect 22465 3547 22523 3553
rect 23566 3544 23572 3596
rect 23624 3584 23630 3596
rect 23860 3584 23888 3615
rect 29822 3612 29828 3624
rect 29880 3612 29886 3664
rect 30558 3612 30564 3664
rect 30616 3652 30622 3664
rect 30926 3652 30932 3664
rect 30616 3624 30932 3652
rect 30616 3612 30622 3624
rect 30926 3612 30932 3624
rect 30984 3612 30990 3664
rect 32861 3655 32919 3661
rect 32861 3621 32873 3655
rect 32907 3621 32919 3655
rect 32861 3615 32919 3621
rect 35253 3655 35311 3661
rect 35253 3621 35265 3655
rect 35299 3621 35311 3655
rect 35253 3615 35311 3621
rect 24581 3587 24639 3593
rect 24581 3584 24593 3587
rect 23624 3556 24593 3584
rect 23624 3544 23630 3556
rect 24581 3553 24593 3556
rect 24627 3553 24639 3587
rect 24581 3547 24639 3553
rect 24946 3544 24952 3596
rect 25004 3584 25010 3596
rect 25869 3587 25927 3593
rect 25869 3584 25881 3587
rect 25004 3556 25881 3584
rect 25004 3544 25010 3556
rect 25869 3553 25881 3556
rect 25915 3553 25927 3587
rect 25869 3547 25927 3553
rect 26145 3587 26203 3593
rect 26145 3553 26157 3587
rect 26191 3584 26203 3587
rect 27801 3587 27859 3593
rect 27801 3584 27813 3587
rect 26191 3556 27813 3584
rect 26191 3553 26203 3556
rect 26145 3547 26203 3553
rect 27801 3553 27813 3556
rect 27847 3584 27859 3587
rect 32674 3584 32680 3596
rect 27847 3556 30052 3584
rect 27847 3553 27859 3556
rect 27801 3547 27859 3553
rect 30024 3528 30052 3556
rect 32140 3556 32680 3584
rect 20027 3488 21312 3516
rect 22005 3519 22063 3525
rect 20027 3485 20039 3488
rect 19981 3479 20039 3485
rect 22005 3485 22017 3519
rect 22051 3516 22063 3519
rect 23290 3516 23296 3528
rect 22051 3488 23296 3516
rect 22051 3485 22063 3488
rect 22005 3479 22063 3485
rect 23290 3476 23296 3488
rect 23348 3476 23354 3528
rect 24394 3476 24400 3528
rect 24452 3516 24458 3528
rect 24489 3519 24547 3525
rect 24489 3516 24501 3519
rect 24452 3488 24501 3516
rect 24452 3476 24458 3488
rect 24489 3485 24501 3488
rect 24535 3485 24547 3519
rect 24489 3479 24547 3485
rect 24765 3519 24823 3525
rect 24765 3485 24777 3519
rect 24811 3516 24823 3519
rect 25222 3516 25228 3528
rect 24811 3488 25228 3516
rect 24811 3485 24823 3488
rect 24765 3479 24823 3485
rect 25222 3476 25228 3488
rect 25280 3476 25286 3528
rect 26694 3476 26700 3528
rect 26752 3516 26758 3528
rect 27341 3519 27399 3525
rect 27341 3516 27353 3519
rect 26752 3488 27353 3516
rect 26752 3476 26758 3488
rect 27341 3485 27353 3488
rect 27387 3485 27399 3519
rect 27982 3516 27988 3528
rect 27943 3488 27988 3516
rect 27341 3479 27399 3485
rect 27982 3476 27988 3488
rect 28040 3476 28046 3528
rect 28169 3519 28227 3525
rect 28169 3485 28181 3519
rect 28215 3516 28227 3519
rect 28813 3519 28871 3525
rect 28813 3516 28825 3519
rect 28215 3488 28825 3516
rect 28215 3485 28227 3488
rect 28169 3479 28227 3485
rect 28813 3485 28825 3488
rect 28859 3485 28871 3519
rect 30006 3516 30012 3528
rect 29967 3488 30012 3516
rect 28813 3479 28871 3485
rect 30006 3476 30012 3488
rect 30064 3476 30070 3528
rect 30101 3519 30159 3525
rect 30101 3485 30113 3519
rect 30147 3516 30159 3519
rect 30190 3516 30196 3528
rect 30147 3488 30196 3516
rect 30147 3485 30159 3488
rect 30101 3479 30159 3485
rect 30190 3476 30196 3488
rect 30248 3476 30254 3528
rect 30745 3519 30803 3525
rect 30745 3485 30757 3519
rect 30791 3516 30803 3519
rect 31018 3516 31024 3528
rect 30791 3488 31024 3516
rect 30791 3485 30803 3488
rect 30745 3479 30803 3485
rect 31018 3476 31024 3488
rect 31076 3476 31082 3528
rect 31846 3516 31852 3528
rect 31807 3488 31852 3516
rect 31846 3476 31852 3488
rect 31904 3476 31910 3528
rect 32030 3516 32036 3528
rect 31991 3488 32036 3516
rect 32030 3476 32036 3488
rect 32088 3476 32094 3528
rect 32140 3525 32168 3556
rect 32674 3544 32680 3556
rect 32732 3544 32738 3596
rect 32876 3528 32904 3615
rect 35268 3584 35296 3615
rect 33980 3556 35296 3584
rect 32125 3519 32183 3525
rect 32125 3485 32137 3519
rect 32171 3485 32183 3519
rect 32125 3479 32183 3485
rect 32214 3476 32220 3528
rect 32272 3516 32278 3528
rect 32272 3488 32317 3516
rect 32272 3476 32278 3488
rect 32858 3476 32864 3528
rect 32916 3476 32922 3528
rect 33042 3516 33048 3528
rect 33003 3488 33048 3516
rect 33042 3476 33048 3488
rect 33100 3476 33106 3528
rect 33778 3516 33784 3528
rect 33691 3488 33784 3516
rect 33778 3476 33784 3488
rect 33836 3476 33842 3528
rect 33980 3525 34008 3556
rect 33965 3519 34023 3525
rect 33965 3485 33977 3519
rect 34011 3485 34023 3519
rect 33965 3479 34023 3485
rect 34422 3476 34428 3528
rect 34480 3516 34486 3528
rect 34698 3516 34704 3528
rect 34480 3488 34704 3516
rect 34480 3476 34486 3488
rect 34698 3476 34704 3488
rect 34756 3476 34762 3528
rect 34790 3476 34796 3528
rect 34848 3516 34854 3528
rect 34977 3519 35035 3525
rect 34977 3516 34989 3519
rect 34848 3488 34989 3516
rect 34848 3476 34854 3488
rect 34977 3485 34989 3488
rect 35023 3485 35035 3519
rect 34977 3479 35035 3485
rect 35069 3519 35127 3525
rect 35069 3485 35081 3519
rect 35115 3516 35127 3519
rect 35434 3516 35440 3528
rect 35115 3488 35440 3516
rect 35115 3485 35127 3488
rect 35069 3479 35127 3485
rect 35434 3476 35440 3488
rect 35492 3476 35498 3528
rect 35710 3516 35716 3528
rect 35671 3488 35716 3516
rect 35710 3476 35716 3488
rect 35768 3476 35774 3528
rect 36538 3516 36544 3528
rect 36499 3488 36544 3516
rect 36538 3476 36544 3488
rect 36596 3476 36602 3528
rect 19337 3451 19395 3457
rect 19337 3417 19349 3451
rect 19383 3448 19395 3451
rect 19518 3448 19524 3460
rect 19383 3420 19524 3448
rect 19383 3417 19395 3420
rect 19337 3411 19395 3417
rect 19518 3408 19524 3420
rect 19576 3408 19582 3460
rect 20248 3451 20306 3457
rect 20248 3417 20260 3451
rect 20294 3448 20306 3451
rect 20898 3448 20904 3460
rect 20294 3420 20904 3448
rect 20294 3417 20306 3420
rect 20248 3411 20306 3417
rect 20898 3408 20904 3420
rect 20956 3408 20962 3460
rect 22710 3451 22768 3457
rect 22710 3448 22722 3451
rect 22066 3420 22722 3448
rect 18322 3380 18328 3392
rect 15896 3352 17540 3380
rect 18283 3352 18328 3380
rect 15896 3340 15902 3352
rect 18322 3340 18328 3352
rect 18380 3340 18386 3392
rect 19242 3340 19248 3392
rect 19300 3380 19306 3392
rect 19429 3383 19487 3389
rect 19429 3380 19441 3383
rect 19300 3352 19441 3380
rect 19300 3340 19306 3352
rect 19429 3349 19441 3352
rect 19475 3349 19487 3383
rect 19429 3343 19487 3349
rect 21821 3383 21879 3389
rect 21821 3349 21833 3383
rect 21867 3380 21879 3383
rect 22066 3380 22094 3420
rect 22710 3417 22722 3420
rect 22756 3417 22768 3451
rect 22710 3411 22768 3417
rect 29822 3408 29828 3460
rect 29880 3448 29886 3460
rect 29880 3420 30972 3448
rect 29880 3408 29886 3420
rect 28626 3380 28632 3392
rect 21867 3352 22094 3380
rect 28587 3352 28632 3380
rect 21867 3349 21879 3352
rect 21821 3343 21879 3349
rect 28626 3340 28632 3352
rect 28684 3340 28690 3392
rect 30285 3383 30343 3389
rect 30285 3349 30297 3383
rect 30331 3380 30343 3383
rect 30834 3380 30840 3392
rect 30331 3352 30840 3380
rect 30331 3349 30343 3352
rect 30285 3343 30343 3349
rect 30834 3340 30840 3352
rect 30892 3340 30898 3392
rect 30944 3389 30972 3420
rect 32950 3408 32956 3460
rect 33008 3448 33014 3460
rect 33796 3448 33824 3476
rect 33008 3420 33824 3448
rect 33008 3408 33014 3420
rect 34330 3408 34336 3460
rect 34388 3448 34394 3460
rect 34885 3451 34943 3457
rect 34885 3448 34897 3451
rect 34388 3420 34897 3448
rect 34388 3408 34394 3420
rect 34885 3417 34897 3420
rect 34931 3417 34943 3451
rect 34885 3411 34943 3417
rect 35158 3408 35164 3460
rect 35216 3448 35222 3460
rect 37921 3451 37979 3457
rect 35216 3420 36860 3448
rect 35216 3408 35222 3420
rect 30929 3383 30987 3389
rect 30929 3349 30941 3383
rect 30975 3349 30987 3383
rect 30929 3343 30987 3349
rect 31110 3340 31116 3392
rect 31168 3380 31174 3392
rect 32214 3380 32220 3392
rect 31168 3352 32220 3380
rect 31168 3340 31174 3352
rect 32214 3340 32220 3352
rect 32272 3340 32278 3392
rect 32306 3340 32312 3392
rect 32364 3380 32370 3392
rect 32401 3383 32459 3389
rect 32401 3380 32413 3383
rect 32364 3352 32413 3380
rect 32364 3340 32370 3352
rect 32401 3349 32413 3352
rect 32447 3349 32459 3383
rect 32401 3343 32459 3349
rect 34149 3383 34207 3389
rect 34149 3349 34161 3383
rect 34195 3380 34207 3383
rect 35250 3380 35256 3392
rect 34195 3352 35256 3380
rect 34195 3349 34207 3352
rect 34149 3343 34207 3349
rect 35250 3340 35256 3352
rect 35308 3340 35314 3392
rect 35434 3340 35440 3392
rect 35492 3380 35498 3392
rect 35897 3383 35955 3389
rect 35897 3380 35909 3383
rect 35492 3352 35909 3380
rect 35492 3340 35498 3352
rect 35897 3349 35909 3352
rect 35943 3349 35955 3383
rect 35897 3343 35955 3349
rect 36446 3340 36452 3392
rect 36504 3380 36510 3392
rect 36725 3383 36783 3389
rect 36725 3380 36737 3383
rect 36504 3352 36737 3380
rect 36504 3340 36510 3352
rect 36725 3349 36737 3352
rect 36771 3349 36783 3383
rect 36832 3380 36860 3420
rect 37921 3417 37933 3451
rect 37967 3448 37979 3451
rect 39390 3448 39396 3460
rect 37967 3420 39396 3448
rect 37967 3417 37979 3420
rect 37921 3411 37979 3417
rect 39390 3408 39396 3420
rect 39448 3408 39454 3460
rect 38013 3383 38071 3389
rect 38013 3380 38025 3383
rect 36832 3352 38025 3380
rect 36725 3343 36783 3349
rect 38013 3349 38025 3352
rect 38059 3349 38071 3383
rect 38013 3343 38071 3349
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 3050 3176 3056 3188
rect 3011 3148 3056 3176
rect 3050 3136 3056 3148
rect 3108 3136 3114 3188
rect 3789 3179 3847 3185
rect 3789 3145 3801 3179
rect 3835 3145 3847 3179
rect 4614 3176 4620 3188
rect 4575 3148 4620 3176
rect 3789 3139 3847 3145
rect 2866 3108 2872 3120
rect 2827 3080 2872 3108
rect 2866 3068 2872 3080
rect 2924 3068 2930 3120
rect 3804 3108 3832 3139
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 5169 3179 5227 3185
rect 5169 3145 5181 3179
rect 5215 3176 5227 3179
rect 5350 3176 5356 3188
rect 5215 3148 5356 3176
rect 5215 3145 5227 3148
rect 5169 3139 5227 3145
rect 5350 3136 5356 3148
rect 5408 3136 5414 3188
rect 6365 3179 6423 3185
rect 6365 3145 6377 3179
rect 6411 3176 6423 3179
rect 8941 3179 8999 3185
rect 6411 3148 8892 3176
rect 6411 3145 6423 3148
rect 6365 3139 6423 3145
rect 3804 3080 5304 3108
rect 1394 3040 1400 3052
rect 1355 3012 1400 3040
rect 1394 3000 1400 3012
rect 1452 3000 1458 3052
rect 3142 3000 3148 3052
rect 3200 3040 3206 3052
rect 3973 3043 4031 3049
rect 3973 3040 3985 3043
rect 3200 3012 3985 3040
rect 3200 3000 3206 3012
rect 3973 3009 3985 3012
rect 4019 3009 4031 3043
rect 3973 3003 4031 3009
rect 4614 3000 4620 3052
rect 4672 3040 4678 3052
rect 4801 3043 4859 3049
rect 4801 3040 4813 3043
rect 4672 3012 4813 3040
rect 4672 3000 4678 3012
rect 4801 3009 4813 3012
rect 4847 3009 4859 3043
rect 4801 3003 4859 3009
rect 5276 2972 5304 3080
rect 5368 3040 5396 3136
rect 8754 3108 8760 3120
rect 7576 3080 8760 3108
rect 5445 3043 5503 3049
rect 5445 3040 5457 3043
rect 5368 3012 5457 3040
rect 5445 3009 5457 3012
rect 5491 3009 5503 3043
rect 5445 3003 5503 3009
rect 6086 3000 6092 3052
rect 6144 3040 6150 3052
rect 7576 3049 7604 3080
rect 8754 3068 8760 3080
rect 8812 3068 8818 3120
rect 6549 3043 6607 3049
rect 6549 3040 6561 3043
rect 6144 3012 6561 3040
rect 6144 3000 6150 3012
rect 6549 3009 6561 3012
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3009 7619 3043
rect 7561 3003 7619 3009
rect 7828 3043 7886 3049
rect 7828 3009 7840 3043
rect 7874 3040 7886 3043
rect 8294 3040 8300 3052
rect 7874 3012 8300 3040
rect 7874 3009 7886 3012
rect 7828 3003 7886 3009
rect 8294 3000 8300 3012
rect 8352 3000 8358 3052
rect 8864 3040 8892 3148
rect 8941 3145 8953 3179
rect 8987 3176 8999 3179
rect 9122 3176 9128 3188
rect 8987 3148 9128 3176
rect 8987 3145 8999 3148
rect 8941 3139 8999 3145
rect 9122 3136 9128 3148
rect 9180 3136 9186 3188
rect 9674 3136 9680 3188
rect 9732 3176 9738 3188
rect 9953 3179 10011 3185
rect 9953 3176 9965 3179
rect 9732 3148 9965 3176
rect 9732 3136 9738 3148
rect 9953 3145 9965 3148
rect 9999 3145 10011 3179
rect 12342 3176 12348 3188
rect 9953 3139 10011 3145
rect 10336 3148 12348 3176
rect 10336 3108 10364 3148
rect 12342 3136 12348 3148
rect 12400 3136 12406 3188
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 12897 3179 12955 3185
rect 12897 3176 12909 3179
rect 12492 3148 12909 3176
rect 12492 3136 12498 3148
rect 12897 3145 12909 3148
rect 12943 3145 12955 3179
rect 12897 3139 12955 3145
rect 14274 3136 14280 3188
rect 14332 3176 14338 3188
rect 15473 3179 15531 3185
rect 15473 3176 15485 3179
rect 14332 3148 15485 3176
rect 14332 3136 14338 3148
rect 15473 3145 15485 3148
rect 15519 3145 15531 3179
rect 15473 3139 15531 3145
rect 16868 3148 18920 3176
rect 10965 3111 11023 3117
rect 10965 3108 10977 3111
rect 10060 3080 10364 3108
rect 10612 3080 10977 3108
rect 9950 3040 9956 3052
rect 8864 3012 9956 3040
rect 9950 3000 9956 3012
rect 10008 3000 10014 3052
rect 5534 2972 5540 2984
rect 5276 2944 5540 2972
rect 5534 2932 5540 2944
rect 5592 2932 5598 2984
rect 10060 2972 10088 3080
rect 10137 3043 10195 3049
rect 10137 3009 10149 3043
rect 10183 3040 10195 3043
rect 10612 3040 10640 3080
rect 10965 3077 10977 3080
rect 11011 3077 11023 3111
rect 11698 3108 11704 3120
rect 11659 3080 11704 3108
rect 10965 3071 11023 3077
rect 11698 3068 11704 3080
rect 11756 3068 11762 3120
rect 11790 3068 11796 3120
rect 11848 3108 11854 3120
rect 12986 3108 12992 3120
rect 11848 3080 11893 3108
rect 12406 3080 12992 3108
rect 11848 3068 11854 3080
rect 10183 3012 10640 3040
rect 10781 3043 10839 3049
rect 10183 3009 10195 3012
rect 10137 3003 10195 3009
rect 10781 3009 10793 3043
rect 10827 3009 10839 3043
rect 10781 3003 10839 3009
rect 8588 2944 10088 2972
rect 10597 2975 10655 2981
rect 2222 2864 2228 2916
rect 2280 2904 2286 2916
rect 3237 2907 3295 2913
rect 2280 2876 2774 2904
rect 2280 2864 2286 2876
rect 934 2796 940 2848
rect 992 2836 998 2848
rect 1581 2839 1639 2845
rect 1581 2836 1593 2839
rect 992 2808 1593 2836
rect 992 2796 998 2808
rect 1581 2805 1593 2808
rect 1627 2805 1639 2839
rect 1581 2799 1639 2805
rect 2038 2796 2044 2848
rect 2096 2836 2102 2848
rect 2317 2839 2375 2845
rect 2317 2836 2329 2839
rect 2096 2808 2329 2836
rect 2096 2796 2102 2808
rect 2317 2805 2329 2808
rect 2363 2805 2375 2839
rect 2746 2836 2774 2876
rect 3237 2873 3249 2907
rect 3283 2904 3295 2907
rect 3283 2876 7604 2904
rect 3283 2873 3295 2876
rect 3237 2867 3295 2873
rect 3053 2839 3111 2845
rect 3053 2836 3065 2839
rect 2746 2808 3065 2836
rect 2317 2799 2375 2805
rect 3053 2805 3065 2808
rect 3099 2805 3111 2839
rect 3053 2799 3111 2805
rect 5350 2796 5356 2848
rect 5408 2836 5414 2848
rect 5629 2839 5687 2845
rect 5629 2836 5641 2839
rect 5408 2808 5641 2836
rect 5408 2796 5414 2808
rect 5629 2805 5641 2808
rect 5675 2805 5687 2839
rect 7576 2836 7604 2876
rect 8588 2836 8616 2944
rect 10597 2941 10609 2975
rect 10643 2972 10655 2975
rect 10796 2972 10824 3003
rect 11146 3000 11152 3052
rect 11204 3040 11210 3052
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 11204 3012 11529 3040
rect 11204 3000 11210 3012
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 11882 3040 11888 3052
rect 11843 3012 11888 3040
rect 11517 3003 11575 3009
rect 11882 3000 11888 3012
rect 11940 3000 11946 3052
rect 12406 3040 12434 3080
rect 12544 3049 12572 3080
rect 12986 3068 12992 3080
rect 13044 3068 13050 3120
rect 13354 3068 13360 3120
rect 13412 3108 13418 3120
rect 13694 3111 13752 3117
rect 13694 3108 13706 3111
rect 13412 3080 13706 3108
rect 13412 3068 13418 3080
rect 13694 3077 13706 3080
rect 13740 3077 13752 3111
rect 13694 3071 13752 3077
rect 14458 3068 14464 3120
rect 14516 3108 14522 3120
rect 16868 3108 16896 3148
rect 14516 3080 16896 3108
rect 14516 3068 14522 3080
rect 12268 3012 12434 3040
rect 12529 3043 12587 3049
rect 10643 2944 10732 2972
rect 10796 2944 12112 2972
rect 10643 2941 10655 2944
rect 10597 2935 10655 2941
rect 9674 2864 9680 2916
rect 9732 2904 9738 2916
rect 10226 2904 10232 2916
rect 9732 2876 10232 2904
rect 9732 2864 9738 2876
rect 10226 2864 10232 2876
rect 10284 2864 10290 2916
rect 10704 2904 10732 2944
rect 12084 2913 12112 2944
rect 12069 2907 12127 2913
rect 10704 2876 10824 2904
rect 7576 2808 8616 2836
rect 5629 2799 5687 2805
rect 9858 2796 9864 2848
rect 9916 2836 9922 2848
rect 10594 2836 10600 2848
rect 9916 2808 10600 2836
rect 9916 2796 9922 2808
rect 10594 2796 10600 2808
rect 10652 2796 10658 2848
rect 10796 2836 10824 2876
rect 12069 2873 12081 2907
rect 12115 2873 12127 2907
rect 12069 2867 12127 2873
rect 12268 2836 12296 3012
rect 12529 3009 12541 3043
rect 12575 3009 12587 3043
rect 12710 3040 12716 3052
rect 12671 3012 12716 3040
rect 12529 3003 12587 3009
rect 12710 3000 12716 3012
rect 12768 3000 12774 3052
rect 13449 3043 13507 3049
rect 13449 3009 13461 3043
rect 13495 3040 13507 3043
rect 13538 3040 13544 3052
rect 13495 3012 13544 3040
rect 13495 3009 13507 3012
rect 13449 3003 13507 3009
rect 13538 3000 13544 3012
rect 13596 3000 13602 3052
rect 15194 3000 15200 3052
rect 15252 3040 15258 3052
rect 15289 3043 15347 3049
rect 15289 3040 15301 3043
rect 15252 3012 15301 3040
rect 15252 3000 15258 3012
rect 15289 3009 15301 3012
rect 15335 3009 15347 3043
rect 15289 3003 15347 3009
rect 16669 3043 16727 3049
rect 16669 3009 16681 3043
rect 16715 3040 16727 3043
rect 16758 3040 16764 3052
rect 16715 3012 16764 3040
rect 16715 3009 16727 3012
rect 16669 3003 16727 3009
rect 16758 3000 16764 3012
rect 16816 3000 16822 3052
rect 16868 3049 16896 3080
rect 16945 3111 17003 3117
rect 16945 3077 16957 3111
rect 16991 3108 17003 3111
rect 17678 3108 17684 3120
rect 16991 3080 17684 3108
rect 16991 3077 17003 3080
rect 16945 3071 17003 3077
rect 17678 3068 17684 3080
rect 17736 3068 17742 3120
rect 18132 3111 18190 3117
rect 18132 3077 18144 3111
rect 18178 3108 18190 3111
rect 18322 3108 18328 3120
rect 18178 3080 18328 3108
rect 18178 3077 18190 3080
rect 18132 3071 18190 3077
rect 18322 3068 18328 3080
rect 18380 3068 18386 3120
rect 16853 3043 16911 3049
rect 16853 3009 16865 3043
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3009 17095 3043
rect 17862 3040 17868 3052
rect 17823 3012 17868 3040
rect 17037 3003 17095 3009
rect 12342 2932 12348 2984
rect 12400 2972 12406 2984
rect 13262 2972 13268 2984
rect 12400 2944 13268 2972
rect 12400 2932 12406 2944
rect 13262 2932 13268 2944
rect 13320 2932 13326 2984
rect 14829 2907 14887 2913
rect 14829 2873 14841 2907
rect 14875 2904 14887 2907
rect 14918 2904 14924 2916
rect 14875 2876 14924 2904
rect 14875 2873 14887 2876
rect 14829 2867 14887 2873
rect 14918 2864 14924 2876
rect 14976 2864 14982 2916
rect 17052 2904 17080 3003
rect 17862 3000 17868 3012
rect 17920 3000 17926 3052
rect 18892 2972 18920 3148
rect 19150 3136 19156 3188
rect 19208 3176 19214 3188
rect 19245 3179 19303 3185
rect 19245 3176 19257 3179
rect 19208 3148 19257 3176
rect 19208 3136 19214 3148
rect 19245 3145 19257 3148
rect 19291 3145 19303 3179
rect 19245 3139 19303 3145
rect 19260 3040 19288 3139
rect 22462 3136 22468 3188
rect 22520 3176 22526 3188
rect 22925 3179 22983 3185
rect 22925 3176 22937 3179
rect 22520 3148 22937 3176
rect 22520 3136 22526 3148
rect 22925 3145 22937 3148
rect 22971 3145 22983 3179
rect 24946 3176 24952 3188
rect 22925 3139 22983 3145
rect 23676 3148 24952 3176
rect 19978 3108 19984 3120
rect 19939 3080 19984 3108
rect 19978 3068 19984 3080
rect 20036 3068 20042 3120
rect 20901 3111 20959 3117
rect 20901 3077 20913 3111
rect 20947 3108 20959 3111
rect 20947 3080 23244 3108
rect 20947 3077 20959 3080
rect 20901 3071 20959 3077
rect 19705 3043 19763 3049
rect 19705 3040 19717 3043
rect 19260 3012 19717 3040
rect 19705 3009 19717 3012
rect 19751 3009 19763 3043
rect 19705 3003 19763 3009
rect 19889 3043 19947 3049
rect 19889 3009 19901 3043
rect 19935 3009 19947 3043
rect 19889 3003 19947 3009
rect 20073 3043 20131 3049
rect 20073 3009 20085 3043
rect 20119 3009 20131 3043
rect 20714 3040 20720 3052
rect 20675 3012 20720 3040
rect 20073 3003 20131 3009
rect 19242 2972 19248 2984
rect 18892 2944 19248 2972
rect 19242 2932 19248 2944
rect 19300 2972 19306 2984
rect 19904 2972 19932 3003
rect 19300 2944 19932 2972
rect 20088 2972 20116 3003
rect 20714 3000 20720 3012
rect 20772 3000 20778 3052
rect 20990 3040 20996 3052
rect 20951 3012 20996 3040
rect 20990 3000 20996 3012
rect 21048 3000 21054 3052
rect 21085 3043 21143 3049
rect 21085 3009 21097 3043
rect 21131 3009 21143 3043
rect 22281 3043 22339 3049
rect 22281 3040 22293 3043
rect 21085 3003 21143 3009
rect 22066 3012 22293 3040
rect 20346 2972 20352 2984
rect 20088 2944 20352 2972
rect 19300 2932 19306 2944
rect 20088 2904 20116 2944
rect 20346 2932 20352 2944
rect 20404 2972 20410 2984
rect 21100 2972 21128 3003
rect 20404 2944 21128 2972
rect 20404 2932 20410 2944
rect 16776 2876 17908 2904
rect 10796 2808 12296 2836
rect 12342 2796 12348 2848
rect 12400 2836 12406 2848
rect 12618 2836 12624 2848
rect 12400 2808 12624 2836
rect 12400 2796 12406 2808
rect 12618 2796 12624 2808
rect 12676 2796 12682 2848
rect 14642 2796 14648 2848
rect 14700 2836 14706 2848
rect 16776 2836 16804 2876
rect 14700 2808 16804 2836
rect 14700 2796 14706 2808
rect 16850 2796 16856 2848
rect 16908 2836 16914 2848
rect 17221 2839 17279 2845
rect 17221 2836 17233 2839
rect 16908 2808 17233 2836
rect 16908 2796 16914 2808
rect 17221 2805 17233 2808
rect 17267 2805 17279 2839
rect 17880 2836 17908 2876
rect 19352 2876 20116 2904
rect 19352 2836 19380 2876
rect 21818 2864 21824 2916
rect 21876 2904 21882 2916
rect 22066 2904 22094 3012
rect 22281 3009 22293 3012
rect 22327 3009 22339 3043
rect 22281 3003 22339 3009
rect 22370 3000 22376 3052
rect 22428 3040 22434 3052
rect 23109 3043 23167 3049
rect 23109 3040 23121 3043
rect 22428 3012 23121 3040
rect 22428 3000 22434 3012
rect 23109 3009 23121 3012
rect 23155 3009 23167 3043
rect 23109 3003 23167 3009
rect 22465 2975 22523 2981
rect 22465 2941 22477 2975
rect 22511 2972 22523 2975
rect 23216 2972 23244 3080
rect 23566 3040 23572 3052
rect 23527 3012 23572 3040
rect 23566 3000 23572 3012
rect 23624 3000 23630 3052
rect 23676 3040 23704 3148
rect 24946 3136 24952 3148
rect 25004 3136 25010 3188
rect 25222 3136 25228 3188
rect 25280 3176 25286 3188
rect 26421 3179 26479 3185
rect 26421 3176 26433 3179
rect 25280 3148 26433 3176
rect 25280 3136 25286 3148
rect 26421 3145 26433 3148
rect 26467 3145 26479 3179
rect 26421 3139 26479 3145
rect 27890 3136 27896 3188
rect 27948 3176 27954 3188
rect 28718 3176 28724 3188
rect 27948 3148 28724 3176
rect 27948 3136 27954 3148
rect 28718 3136 28724 3148
rect 28776 3136 28782 3188
rect 28810 3136 28816 3188
rect 28868 3176 28874 3188
rect 35158 3176 35164 3188
rect 28868 3148 35164 3176
rect 28868 3136 28874 3148
rect 35158 3136 35164 3148
rect 35216 3136 35222 3188
rect 36541 3179 36599 3185
rect 36541 3145 36553 3179
rect 36587 3145 36599 3179
rect 36541 3139 36599 3145
rect 23842 3108 23848 3120
rect 23803 3080 23848 3108
rect 23842 3068 23848 3080
rect 23900 3068 23906 3120
rect 27608 3111 27666 3117
rect 25056 3080 27384 3108
rect 25056 3052 25084 3080
rect 23753 3043 23811 3049
rect 23753 3040 23765 3043
rect 23676 3012 23765 3040
rect 23676 2972 23704 3012
rect 23753 3009 23765 3012
rect 23799 3009 23811 3043
rect 23753 3003 23811 3009
rect 23937 3043 23995 3049
rect 23937 3009 23949 3043
rect 23983 3040 23995 3043
rect 24854 3040 24860 3052
rect 23983 3012 24860 3040
rect 23983 3009 23995 3012
rect 23937 3003 23995 3009
rect 22511 2944 23704 2972
rect 22511 2941 22523 2944
rect 22465 2935 22523 2941
rect 21876 2876 22094 2904
rect 21876 2864 21882 2876
rect 17880 2808 19380 2836
rect 17221 2799 17279 2805
rect 19426 2796 19432 2848
rect 19484 2836 19490 2848
rect 20257 2839 20315 2845
rect 20257 2836 20269 2839
rect 19484 2808 20269 2836
rect 19484 2796 19490 2808
rect 20257 2805 20269 2808
rect 20303 2805 20315 2839
rect 20257 2799 20315 2805
rect 20806 2796 20812 2848
rect 20864 2836 20870 2848
rect 21269 2839 21327 2845
rect 21269 2836 21281 2839
rect 20864 2808 21281 2836
rect 20864 2796 20870 2808
rect 21269 2805 21281 2808
rect 21315 2805 21327 2839
rect 21269 2799 21327 2805
rect 23474 2796 23480 2848
rect 23532 2836 23538 2848
rect 24121 2839 24179 2845
rect 24121 2836 24133 2839
rect 23532 2808 24133 2836
rect 23532 2796 23538 2808
rect 24121 2805 24133 2808
rect 24167 2805 24179 2839
rect 24596 2836 24624 3012
rect 24854 3000 24860 3012
rect 24912 3000 24918 3052
rect 25038 3040 25044 3052
rect 24999 3012 25044 3040
rect 25038 3000 25044 3012
rect 25096 3000 25102 3052
rect 25314 3049 25320 3052
rect 25308 3040 25320 3049
rect 25275 3012 25320 3040
rect 25308 3003 25320 3012
rect 25314 3000 25320 3003
rect 25372 3000 25378 3052
rect 27356 3049 27384 3080
rect 27608 3077 27620 3111
rect 27654 3108 27666 3111
rect 28626 3108 28632 3120
rect 27654 3080 28632 3108
rect 27654 3077 27666 3080
rect 27608 3071 27666 3077
rect 28626 3068 28632 3080
rect 28684 3068 28690 3120
rect 30006 3068 30012 3120
rect 30064 3108 30070 3120
rect 32030 3108 32036 3120
rect 30064 3080 32036 3108
rect 30064 3068 30070 3080
rect 32030 3068 32036 3080
rect 32088 3068 32094 3120
rect 34232 3111 34290 3117
rect 32140 3080 34008 3108
rect 27341 3043 27399 3049
rect 27341 3009 27353 3043
rect 27387 3009 27399 3043
rect 29638 3040 29644 3052
rect 29599 3012 29644 3040
rect 27341 3003 27399 3009
rect 29638 3000 29644 3012
rect 29696 3000 29702 3052
rect 29908 3043 29966 3049
rect 29908 3009 29920 3043
rect 29954 3040 29966 3043
rect 30926 3040 30932 3052
rect 29954 3012 30932 3040
rect 29954 3009 29966 3012
rect 29908 3003 29966 3009
rect 30926 3000 30932 3012
rect 30984 3000 30990 3052
rect 31570 3000 31576 3052
rect 31628 3040 31634 3052
rect 32140 3049 32168 3080
rect 32125 3043 32183 3049
rect 32125 3040 32137 3043
rect 31628 3012 32137 3040
rect 31628 3000 31634 3012
rect 32125 3009 32137 3012
rect 32171 3009 32183 3043
rect 32125 3003 32183 3009
rect 32392 3043 32450 3049
rect 32392 3009 32404 3043
rect 32438 3040 32450 3043
rect 32858 3040 32864 3052
rect 32438 3012 32864 3040
rect 32438 3009 32450 3012
rect 32392 3003 32450 3009
rect 32858 3000 32864 3012
rect 32916 3000 32922 3052
rect 33980 3049 34008 3080
rect 34232 3077 34244 3111
rect 34278 3108 34290 3111
rect 36556 3108 36584 3139
rect 34278 3080 35204 3108
rect 34278 3077 34290 3080
rect 34232 3071 34290 3077
rect 33965 3043 34023 3049
rect 33965 3009 33977 3043
rect 34011 3009 34023 3043
rect 35176 3040 35204 3080
rect 35452 3080 36584 3108
rect 35452 3040 35480 3080
rect 35176 3012 35480 3040
rect 33965 3003 34023 3009
rect 35526 3000 35532 3052
rect 35584 3040 35590 3052
rect 35805 3043 35863 3049
rect 35805 3040 35817 3043
rect 35584 3012 35817 3040
rect 35584 3000 35590 3012
rect 35805 3009 35817 3012
rect 35851 3009 35863 3043
rect 35805 3003 35863 3009
rect 36725 3043 36783 3049
rect 36725 3009 36737 3043
rect 36771 3009 36783 3043
rect 36725 3003 36783 3009
rect 37277 3043 37335 3049
rect 37277 3009 37289 3043
rect 37323 3040 37335 3043
rect 38286 3040 38292 3052
rect 37323 3012 38292 3040
rect 37323 3009 37335 3012
rect 37277 3003 37335 3009
rect 35250 2932 35256 2984
rect 35308 2972 35314 2984
rect 36740 2972 36768 3003
rect 38286 3000 38292 3012
rect 38344 3000 38350 3052
rect 35308 2944 36768 2972
rect 35308 2932 35314 2944
rect 36906 2932 36912 2984
rect 36964 2972 36970 2984
rect 37553 2975 37611 2981
rect 37553 2972 37565 2975
rect 36964 2944 37565 2972
rect 36964 2932 36970 2944
rect 37553 2941 37565 2944
rect 37599 2941 37611 2975
rect 37553 2935 37611 2941
rect 31386 2904 31392 2916
rect 30576 2876 31392 2904
rect 25774 2836 25780 2848
rect 24596 2808 25780 2836
rect 24121 2799 24179 2805
rect 25774 2796 25780 2808
rect 25832 2796 25838 2848
rect 28074 2796 28080 2848
rect 28132 2836 28138 2848
rect 30576 2836 30604 2876
rect 31386 2864 31392 2876
rect 31444 2864 31450 2916
rect 31018 2836 31024 2848
rect 28132 2808 30604 2836
rect 30979 2808 31024 2836
rect 28132 2796 28138 2808
rect 31018 2796 31024 2808
rect 31076 2796 31082 2848
rect 31846 2796 31852 2848
rect 31904 2836 31910 2848
rect 33505 2839 33563 2845
rect 33505 2836 33517 2839
rect 31904 2808 33517 2836
rect 31904 2796 31910 2808
rect 33505 2805 33517 2808
rect 33551 2805 33563 2839
rect 33505 2799 33563 2805
rect 34698 2796 34704 2848
rect 34756 2836 34762 2848
rect 35345 2839 35403 2845
rect 35345 2836 35357 2839
rect 34756 2808 35357 2836
rect 34756 2796 34762 2808
rect 35345 2805 35357 2808
rect 35391 2805 35403 2839
rect 35986 2836 35992 2848
rect 35947 2808 35992 2836
rect 35345 2799 35403 2805
rect 35986 2796 35992 2808
rect 36044 2796 36050 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 2639 2635 2697 2641
rect 2639 2601 2651 2635
rect 2685 2632 2697 2635
rect 14826 2632 14832 2644
rect 2685 2604 13124 2632
rect 14787 2604 14832 2632
rect 2685 2601 2697 2604
rect 2639 2595 2697 2601
rect 12158 2564 12164 2576
rect 3988 2536 12164 2564
rect 1946 2496 1952 2508
rect 1907 2468 1952 2496
rect 1946 2456 1952 2468
rect 2004 2456 2010 2508
rect 2409 2499 2467 2505
rect 2409 2465 2421 2499
rect 2455 2496 2467 2499
rect 2774 2496 2780 2508
rect 2455 2468 2780 2496
rect 2455 2465 2467 2468
rect 2409 2459 2467 2465
rect 2774 2456 2780 2468
rect 2832 2456 2838 2508
rect 3988 2437 4016 2536
rect 12158 2524 12164 2536
rect 12216 2524 12222 2576
rect 5258 2496 5264 2508
rect 5219 2468 5264 2496
rect 5258 2456 5264 2468
rect 5316 2456 5322 2508
rect 11422 2496 11428 2508
rect 8772 2468 11428 2496
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2397 4031 2431
rect 4982 2428 4988 2440
rect 4943 2400 4988 2428
rect 3973 2391 4031 2397
rect 4982 2388 4988 2400
rect 5040 2388 5046 2440
rect 6914 2388 6920 2440
rect 6972 2428 6978 2440
rect 6972 2400 7017 2428
rect 6972 2388 6978 2400
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 7837 2431 7895 2437
rect 7837 2428 7849 2431
rect 7616 2400 7849 2428
rect 7616 2388 7622 2400
rect 7837 2397 7849 2400
rect 7883 2397 7895 2431
rect 7837 2391 7895 2397
rect 566 2320 572 2372
rect 624 2360 630 2372
rect 1765 2363 1823 2369
rect 1765 2360 1777 2363
rect 624 2332 1777 2360
rect 624 2320 630 2332
rect 1765 2329 1777 2332
rect 1811 2329 1823 2363
rect 8772 2360 8800 2468
rect 11422 2456 11428 2468
rect 11480 2456 11486 2508
rect 8938 2428 8944 2440
rect 8899 2400 8944 2428
rect 8938 2388 8944 2400
rect 8996 2388 9002 2440
rect 9861 2431 9919 2437
rect 9861 2397 9873 2431
rect 9907 2428 9919 2431
rect 10318 2428 10324 2440
rect 9907 2400 10324 2428
rect 9907 2397 9919 2400
rect 9861 2391 9919 2397
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 10781 2431 10839 2437
rect 10781 2397 10793 2431
rect 10827 2397 10839 2431
rect 11514 2428 11520 2440
rect 11475 2400 11520 2428
rect 10781 2391 10839 2397
rect 1765 2323 1823 2329
rect 7668 2332 8800 2360
rect 3878 2252 3884 2304
rect 3936 2292 3942 2304
rect 4157 2295 4215 2301
rect 4157 2292 4169 2295
rect 3936 2264 4169 2292
rect 3936 2252 3942 2264
rect 4157 2261 4169 2264
rect 4203 2261 4215 2295
rect 4157 2255 4215 2261
rect 6822 2252 6828 2304
rect 6880 2292 6886 2304
rect 7668 2301 7696 2332
rect 9030 2320 9036 2372
rect 9088 2360 9094 2372
rect 10796 2360 10824 2391
rect 11514 2388 11520 2400
rect 11572 2388 11578 2440
rect 12253 2431 12311 2437
rect 12253 2397 12265 2431
rect 12299 2428 12311 2431
rect 12986 2428 12992 2440
rect 12299 2400 12992 2428
rect 12299 2397 12311 2400
rect 12253 2391 12311 2397
rect 12986 2388 12992 2400
rect 13044 2388 13050 2440
rect 9088 2332 10824 2360
rect 13096 2360 13124 2604
rect 14826 2592 14832 2604
rect 14884 2592 14890 2644
rect 17034 2632 17040 2644
rect 16995 2604 17040 2632
rect 17034 2592 17040 2604
rect 17092 2592 17098 2644
rect 19518 2592 19524 2644
rect 19576 2632 19582 2644
rect 19613 2635 19671 2641
rect 19613 2632 19625 2635
rect 19576 2604 19625 2632
rect 19576 2592 19582 2604
rect 19613 2601 19625 2604
rect 19659 2601 19671 2635
rect 19613 2595 19671 2601
rect 20993 2635 21051 2641
rect 20993 2601 21005 2635
rect 21039 2632 21051 2635
rect 21082 2632 21088 2644
rect 21039 2604 21088 2632
rect 21039 2601 21051 2604
rect 20993 2595 21051 2601
rect 21082 2592 21088 2604
rect 21140 2592 21146 2644
rect 23290 2592 23296 2644
rect 23348 2632 23354 2644
rect 23661 2635 23719 2641
rect 23661 2632 23673 2635
rect 23348 2604 23673 2632
rect 23348 2592 23354 2604
rect 23661 2601 23673 2604
rect 23707 2601 23719 2635
rect 23661 2595 23719 2601
rect 24857 2635 24915 2641
rect 24857 2601 24869 2635
rect 24903 2632 24915 2635
rect 25590 2632 25596 2644
rect 24903 2604 25596 2632
rect 24903 2601 24915 2604
rect 24857 2595 24915 2601
rect 25590 2592 25596 2604
rect 25648 2592 25654 2644
rect 25700 2604 27016 2632
rect 18874 2564 18880 2576
rect 15856 2536 18880 2564
rect 14918 2496 14924 2508
rect 14292 2468 14924 2496
rect 13173 2431 13231 2437
rect 13173 2397 13185 2431
rect 13219 2428 13231 2431
rect 14182 2428 14188 2440
rect 13219 2400 14188 2428
rect 13219 2397 13231 2400
rect 13173 2391 13231 2397
rect 14182 2388 14188 2400
rect 14240 2388 14246 2440
rect 14292 2437 14320 2468
rect 14918 2456 14924 2468
rect 14976 2456 14982 2508
rect 14277 2431 14335 2437
rect 14277 2397 14289 2431
rect 14323 2397 14335 2431
rect 14458 2428 14464 2440
rect 14419 2400 14464 2428
rect 14277 2391 14335 2397
rect 14458 2388 14464 2400
rect 14516 2388 14522 2440
rect 14642 2428 14648 2440
rect 14603 2400 14648 2428
rect 14642 2388 14648 2400
rect 14700 2388 14706 2440
rect 15856 2437 15884 2536
rect 18874 2524 18880 2536
rect 18932 2524 18938 2576
rect 20898 2524 20904 2576
rect 20956 2564 20962 2576
rect 22741 2567 22799 2573
rect 22741 2564 22753 2567
rect 20956 2536 22753 2564
rect 20956 2524 20962 2536
rect 22741 2533 22753 2536
rect 22787 2533 22799 2567
rect 22741 2527 22799 2533
rect 24302 2524 24308 2576
rect 24360 2564 24366 2576
rect 25700 2564 25728 2604
rect 24360 2536 25728 2564
rect 25869 2567 25927 2573
rect 24360 2524 24366 2536
rect 25869 2533 25881 2567
rect 25915 2533 25927 2567
rect 25869 2527 25927 2533
rect 16669 2499 16727 2505
rect 16669 2465 16681 2499
rect 16715 2496 16727 2499
rect 19245 2499 19303 2505
rect 19245 2496 19257 2499
rect 16715 2468 19257 2496
rect 16715 2465 16727 2468
rect 16669 2459 16727 2465
rect 19245 2465 19257 2468
rect 19291 2496 19303 2499
rect 20625 2499 20683 2505
rect 20625 2496 20637 2499
rect 19291 2468 20637 2496
rect 19291 2465 19303 2468
rect 19245 2459 19303 2465
rect 20625 2465 20637 2468
rect 20671 2496 20683 2499
rect 23293 2499 23351 2505
rect 23293 2496 23305 2499
rect 20671 2468 23305 2496
rect 20671 2465 20683 2468
rect 20625 2459 20683 2465
rect 23293 2465 23305 2468
rect 23339 2496 23351 2499
rect 24486 2496 24492 2508
rect 23339 2468 24492 2496
rect 23339 2465 23351 2468
rect 23293 2459 23351 2465
rect 24486 2456 24492 2468
rect 24544 2456 24550 2508
rect 25884 2496 25912 2527
rect 24688 2468 25912 2496
rect 15841 2431 15899 2437
rect 15841 2397 15853 2431
rect 15887 2397 15899 2431
rect 16850 2428 16856 2440
rect 16811 2400 16856 2428
rect 15841 2391 15899 2397
rect 16850 2388 16856 2400
rect 16908 2388 16914 2440
rect 17681 2431 17739 2437
rect 17681 2397 17693 2431
rect 17727 2428 17739 2431
rect 18230 2428 18236 2440
rect 17727 2400 18236 2428
rect 17727 2397 17739 2400
rect 17681 2391 17739 2397
rect 18230 2388 18236 2400
rect 18288 2388 18294 2440
rect 18417 2431 18475 2437
rect 18417 2397 18429 2431
rect 18463 2397 18475 2431
rect 19426 2428 19432 2440
rect 19387 2400 19432 2428
rect 18417 2391 18475 2397
rect 14553 2363 14611 2369
rect 13096 2332 13492 2360
rect 9088 2320 9094 2332
rect 7101 2295 7159 2301
rect 7101 2292 7113 2295
rect 6880 2264 7113 2292
rect 6880 2252 6886 2264
rect 7101 2261 7113 2264
rect 7147 2261 7159 2295
rect 7101 2255 7159 2261
rect 7653 2295 7711 2301
rect 7653 2261 7665 2295
rect 7699 2261 7711 2295
rect 7653 2255 7711 2261
rect 8294 2252 8300 2304
rect 8352 2292 8358 2304
rect 9125 2295 9183 2301
rect 9125 2292 9137 2295
rect 8352 2264 9137 2292
rect 8352 2252 8358 2264
rect 9125 2261 9137 2264
rect 9171 2261 9183 2295
rect 9125 2255 9183 2261
rect 9766 2252 9772 2304
rect 9824 2292 9830 2304
rect 10045 2295 10103 2301
rect 10045 2292 10057 2295
rect 9824 2264 10057 2292
rect 9824 2252 9830 2264
rect 10045 2261 10057 2264
rect 10091 2261 10103 2295
rect 10594 2292 10600 2304
rect 10555 2264 10600 2292
rect 10045 2255 10103 2261
rect 10594 2252 10600 2264
rect 10652 2252 10658 2304
rect 10870 2252 10876 2304
rect 10928 2292 10934 2304
rect 11701 2295 11759 2301
rect 11701 2292 11713 2295
rect 10928 2264 11713 2292
rect 10928 2252 10934 2264
rect 11701 2261 11713 2264
rect 11747 2261 11759 2295
rect 11701 2255 11759 2261
rect 11974 2252 11980 2304
rect 12032 2292 12038 2304
rect 12437 2295 12495 2301
rect 12437 2292 12449 2295
rect 12032 2264 12449 2292
rect 12032 2252 12038 2264
rect 12437 2261 12449 2264
rect 12483 2261 12495 2295
rect 12437 2255 12495 2261
rect 13078 2252 13084 2304
rect 13136 2292 13142 2304
rect 13357 2295 13415 2301
rect 13357 2292 13369 2295
rect 13136 2264 13369 2292
rect 13136 2252 13142 2264
rect 13357 2261 13369 2264
rect 13403 2261 13415 2295
rect 13464 2292 13492 2332
rect 14553 2329 14565 2363
rect 14599 2360 14611 2363
rect 15746 2360 15752 2372
rect 14599 2332 15752 2360
rect 14599 2329 14611 2332
rect 14553 2323 14611 2329
rect 15746 2320 15752 2332
rect 15804 2320 15810 2372
rect 18138 2360 18144 2372
rect 15856 2332 18144 2360
rect 15856 2292 15884 2332
rect 18138 2320 18144 2332
rect 18196 2320 18202 2372
rect 18432 2360 18460 2391
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 20806 2428 20812 2440
rect 20767 2400 20812 2428
rect 20806 2388 20812 2400
rect 20864 2388 20870 2440
rect 21821 2431 21879 2437
rect 21821 2428 21833 2431
rect 20916 2400 21833 2428
rect 20254 2360 20260 2372
rect 18432 2332 20260 2360
rect 20254 2320 20260 2332
rect 20312 2320 20318 2372
rect 20438 2320 20444 2372
rect 20496 2360 20502 2372
rect 20916 2360 20944 2400
rect 21821 2397 21833 2400
rect 21867 2397 21879 2431
rect 22557 2431 22615 2437
rect 22557 2428 22569 2431
rect 21821 2391 21879 2397
rect 22066 2400 22569 2428
rect 20496 2332 20944 2360
rect 20496 2320 20502 2332
rect 21174 2320 21180 2372
rect 21232 2360 21238 2372
rect 22066 2360 22094 2400
rect 22557 2397 22569 2400
rect 22603 2397 22615 2431
rect 23474 2428 23480 2440
rect 23435 2400 23480 2428
rect 22557 2391 22615 2397
rect 23474 2388 23480 2400
rect 23532 2388 23538 2440
rect 24688 2437 24716 2468
rect 24673 2431 24731 2437
rect 24673 2397 24685 2431
rect 24719 2397 24731 2431
rect 24673 2391 24731 2397
rect 25222 2388 25228 2440
rect 25280 2428 25286 2440
rect 25317 2431 25375 2437
rect 25317 2428 25329 2431
rect 25280 2400 25329 2428
rect 25280 2388 25286 2400
rect 25317 2397 25329 2400
rect 25363 2397 25375 2431
rect 25317 2391 25375 2397
rect 25685 2431 25743 2437
rect 25685 2397 25697 2431
rect 25731 2428 25743 2431
rect 25774 2428 25780 2440
rect 25731 2400 25780 2428
rect 25731 2397 25743 2400
rect 25685 2391 25743 2397
rect 25774 2388 25780 2400
rect 25832 2388 25838 2440
rect 26988 2437 27016 2604
rect 27982 2592 27988 2644
rect 28040 2632 28046 2644
rect 28445 2635 28503 2641
rect 28445 2632 28457 2635
rect 28040 2604 28457 2632
rect 28040 2592 28046 2604
rect 28445 2601 28457 2604
rect 28491 2601 28503 2635
rect 30190 2632 30196 2644
rect 30151 2604 30196 2632
rect 28445 2595 28503 2601
rect 30190 2592 30196 2604
rect 30248 2592 30254 2644
rect 30926 2592 30932 2644
rect 30984 2632 30990 2644
rect 31389 2635 31447 2641
rect 31389 2632 31401 2635
rect 30984 2604 31401 2632
rect 30984 2592 30990 2604
rect 31389 2601 31401 2604
rect 31435 2601 31447 2635
rect 31389 2595 31447 2601
rect 32493 2635 32551 2641
rect 32493 2601 32505 2635
rect 32539 2632 32551 2635
rect 33042 2632 33048 2644
rect 32539 2604 33048 2632
rect 32539 2601 32551 2604
rect 32493 2595 32551 2601
rect 33042 2592 33048 2604
rect 33100 2592 33106 2644
rect 30374 2564 30380 2576
rect 28000 2536 29592 2564
rect 28000 2440 28028 2536
rect 26979 2431 27037 2437
rect 26979 2397 26991 2431
rect 27025 2397 27037 2431
rect 27890 2428 27896 2440
rect 27851 2400 27896 2428
rect 26979 2391 27037 2397
rect 27890 2388 27896 2400
rect 27948 2388 27954 2440
rect 27982 2388 27988 2440
rect 28040 2430 28046 2440
rect 28077 2431 28135 2437
rect 28077 2430 28089 2431
rect 28040 2402 28089 2430
rect 28040 2388 28046 2402
rect 28077 2397 28089 2402
rect 28123 2397 28135 2431
rect 28258 2428 28264 2440
rect 28219 2400 28264 2428
rect 28077 2391 28135 2397
rect 28258 2388 28264 2400
rect 28316 2388 28322 2440
rect 21232 2332 22094 2360
rect 21232 2320 21238 2332
rect 24854 2320 24860 2372
rect 24912 2360 24918 2372
rect 25498 2360 25504 2372
rect 24912 2332 25504 2360
rect 24912 2320 24918 2332
rect 25498 2320 25504 2332
rect 25556 2320 25562 2372
rect 25593 2363 25651 2369
rect 25593 2329 25605 2363
rect 25639 2360 25651 2363
rect 27338 2360 27344 2372
rect 25639 2332 27344 2360
rect 25639 2329 25651 2332
rect 25593 2323 25651 2329
rect 27338 2320 27344 2332
rect 27396 2320 27402 2372
rect 28169 2363 28227 2369
rect 28169 2329 28181 2363
rect 28215 2360 28227 2363
rect 29454 2360 29460 2372
rect 28215 2332 29460 2360
rect 28215 2329 28227 2332
rect 28169 2323 28227 2329
rect 29454 2320 29460 2332
rect 29512 2320 29518 2372
rect 29564 2360 29592 2536
rect 29656 2536 30380 2564
rect 29656 2437 29684 2536
rect 30374 2524 30380 2536
rect 30432 2564 30438 2576
rect 31018 2564 31024 2576
rect 30432 2536 31024 2564
rect 30432 2524 30438 2536
rect 31018 2524 31024 2536
rect 31076 2524 31082 2576
rect 32950 2564 32956 2576
rect 32140 2536 32956 2564
rect 31110 2496 31116 2508
rect 30024 2468 31116 2496
rect 30024 2440 30052 2468
rect 31110 2456 31116 2468
rect 31168 2456 31174 2508
rect 32030 2456 32036 2508
rect 32088 2496 32094 2508
rect 32140 2505 32168 2536
rect 32950 2524 32956 2536
rect 33008 2524 33014 2576
rect 33134 2524 33140 2576
rect 33192 2564 33198 2576
rect 34885 2567 34943 2573
rect 34885 2564 34897 2567
rect 33192 2536 34897 2564
rect 33192 2524 33198 2536
rect 34885 2533 34897 2536
rect 34931 2533 34943 2567
rect 34885 2527 34943 2533
rect 32125 2499 32183 2505
rect 32125 2496 32137 2499
rect 32088 2468 32137 2496
rect 32088 2456 32094 2468
rect 32125 2465 32137 2468
rect 32171 2465 32183 2499
rect 32125 2459 32183 2465
rect 32214 2456 32220 2508
rect 32272 2496 32278 2508
rect 32272 2468 32996 2496
rect 32272 2456 32278 2468
rect 29641 2431 29699 2437
rect 29641 2397 29653 2431
rect 29687 2397 29699 2431
rect 30006 2428 30012 2440
rect 29919 2400 30012 2428
rect 29641 2391 29699 2397
rect 30006 2388 30012 2400
rect 30064 2388 30070 2440
rect 30650 2428 30656 2440
rect 30611 2400 30656 2428
rect 30650 2388 30656 2400
rect 30708 2388 30714 2440
rect 30834 2388 30840 2440
rect 30892 2428 30898 2440
rect 31573 2431 31631 2437
rect 31573 2428 31585 2431
rect 30892 2400 31585 2428
rect 30892 2388 30898 2400
rect 31573 2397 31585 2400
rect 31619 2397 31631 2431
rect 32306 2428 32312 2440
rect 32267 2400 32312 2428
rect 31573 2391 31631 2397
rect 32306 2388 32312 2400
rect 32364 2388 32370 2440
rect 32968 2437 32996 2468
rect 33042 2456 33048 2508
rect 33100 2496 33106 2508
rect 37553 2499 37611 2505
rect 37553 2496 37565 2499
rect 33100 2468 37565 2496
rect 33100 2456 33106 2468
rect 37553 2465 37565 2468
rect 37599 2465 37611 2499
rect 37553 2459 37611 2465
rect 32953 2431 33011 2437
rect 32953 2397 32965 2431
rect 32999 2397 33011 2431
rect 33686 2428 33692 2440
rect 33647 2400 33692 2428
rect 32953 2391 33011 2397
rect 33686 2388 33692 2400
rect 33744 2388 33750 2440
rect 33778 2388 33784 2440
rect 33836 2428 33842 2440
rect 34701 2431 34759 2437
rect 34701 2428 34713 2431
rect 33836 2400 34713 2428
rect 33836 2388 33842 2400
rect 34701 2397 34713 2400
rect 34747 2397 34759 2431
rect 34701 2391 34759 2397
rect 35897 2431 35955 2437
rect 35897 2397 35909 2431
rect 35943 2428 35955 2431
rect 36078 2428 36084 2440
rect 35943 2400 36084 2428
rect 35943 2397 35955 2400
rect 35897 2391 35955 2397
rect 36078 2388 36084 2400
rect 36136 2388 36142 2440
rect 36170 2388 36176 2440
rect 36228 2428 36234 2440
rect 36228 2400 36273 2428
rect 36228 2388 36234 2400
rect 37182 2388 37188 2440
rect 37240 2428 37246 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 37240 2400 37289 2428
rect 37240 2388 37246 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 29825 2363 29883 2369
rect 29825 2360 29837 2363
rect 29564 2332 29837 2360
rect 29825 2329 29837 2332
rect 29871 2329 29883 2363
rect 29825 2323 29883 2329
rect 29917 2363 29975 2369
rect 29917 2329 29929 2363
rect 29963 2360 29975 2363
rect 31478 2360 31484 2372
rect 29963 2332 31484 2360
rect 29963 2329 29975 2332
rect 29917 2323 29975 2329
rect 31478 2320 31484 2332
rect 31536 2320 31542 2372
rect 32030 2320 32036 2372
rect 32088 2360 32094 2372
rect 32088 2332 33916 2360
rect 32088 2320 32094 2332
rect 13464 2264 15884 2292
rect 16025 2295 16083 2301
rect 13357 2255 13415 2261
rect 16025 2261 16037 2295
rect 16071 2292 16083 2295
rect 16482 2292 16488 2304
rect 16071 2264 16488 2292
rect 16071 2261 16083 2264
rect 16025 2255 16083 2261
rect 16482 2252 16488 2264
rect 16540 2252 16546 2304
rect 17586 2252 17592 2304
rect 17644 2292 17650 2304
rect 17865 2295 17923 2301
rect 17865 2292 17877 2295
rect 17644 2264 17877 2292
rect 17644 2252 17650 2264
rect 17865 2261 17877 2264
rect 17911 2261 17923 2295
rect 17865 2255 17923 2261
rect 18601 2295 18659 2301
rect 18601 2261 18613 2295
rect 18647 2292 18659 2295
rect 18690 2292 18696 2304
rect 18647 2264 18696 2292
rect 18647 2261 18659 2264
rect 18601 2255 18659 2261
rect 18690 2252 18696 2264
rect 18748 2252 18754 2304
rect 20070 2252 20076 2304
rect 20128 2292 20134 2304
rect 22005 2295 22063 2301
rect 22005 2292 22017 2295
rect 20128 2264 22017 2292
rect 20128 2252 20134 2264
rect 22005 2261 22017 2264
rect 22051 2261 22063 2295
rect 22005 2255 22063 2261
rect 24210 2252 24216 2304
rect 24268 2292 24274 2304
rect 27157 2295 27215 2301
rect 27157 2292 27169 2295
rect 24268 2264 27169 2292
rect 24268 2252 24274 2264
rect 27157 2261 27169 2264
rect 27203 2261 27215 2295
rect 27157 2255 27215 2261
rect 28718 2252 28724 2304
rect 28776 2292 28782 2304
rect 30837 2295 30895 2301
rect 30837 2292 30849 2295
rect 28776 2264 30849 2292
rect 28776 2252 28782 2264
rect 30837 2261 30849 2264
rect 30883 2261 30895 2295
rect 30837 2255 30895 2261
rect 30926 2252 30932 2304
rect 30984 2292 30990 2304
rect 33888 2301 33916 2332
rect 33137 2295 33195 2301
rect 33137 2292 33149 2295
rect 30984 2264 33149 2292
rect 30984 2252 30990 2264
rect 33137 2261 33149 2264
rect 33183 2261 33195 2295
rect 33137 2255 33195 2261
rect 33873 2295 33931 2301
rect 33873 2261 33885 2295
rect 33919 2261 33931 2295
rect 33873 2255 33931 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 6914 2048 6920 2100
rect 6972 2088 6978 2100
rect 10962 2088 10968 2100
rect 6972 2060 10968 2088
rect 6972 2048 6978 2060
rect 10962 2048 10968 2060
rect 11020 2048 11026 2100
rect 11514 2048 11520 2100
rect 11572 2088 11578 2100
rect 16574 2088 16580 2100
rect 11572 2060 16580 2088
rect 11572 2048 11578 2060
rect 16574 2048 16580 2060
rect 16632 2048 16638 2100
rect 25498 2048 25504 2100
rect 25556 2088 25562 2100
rect 27982 2088 27988 2100
rect 25556 2060 27988 2088
rect 25556 2048 25562 2060
rect 27982 2048 27988 2060
rect 28040 2048 28046 2100
rect 28166 2048 28172 2100
rect 28224 2088 28230 2100
rect 33686 2088 33692 2100
rect 28224 2060 33692 2088
rect 28224 2048 28230 2060
rect 33686 2048 33692 2060
rect 33744 2048 33750 2100
rect 8938 1980 8944 2032
rect 8996 2020 9002 2032
rect 15930 2020 15936 2032
rect 8996 1992 15936 2020
rect 8996 1980 9002 1992
rect 15930 1980 15936 1992
rect 15988 1980 15994 2032
rect 26602 1980 26608 2032
rect 26660 2020 26666 2032
rect 33042 2020 33048 2032
rect 26660 1992 33048 2020
rect 26660 1980 26666 1992
rect 33042 1980 33048 1992
rect 33100 1980 33106 2032
rect 25774 1912 25780 1964
rect 25832 1952 25838 1964
rect 28258 1952 28264 1964
rect 25832 1924 28264 1952
rect 25832 1912 25838 1924
rect 28258 1912 28264 1924
rect 28316 1952 28322 1964
rect 30006 1952 30012 1964
rect 28316 1924 30012 1952
rect 28316 1912 28322 1924
rect 30006 1912 30012 1924
rect 30064 1912 30070 1964
rect 24578 1368 24584 1420
rect 24636 1408 24642 1420
rect 27430 1408 27436 1420
rect 24636 1380 27436 1408
rect 24636 1368 24642 1380
rect 27430 1368 27436 1380
rect 27488 1368 27494 1420
rect 34238 1368 34244 1420
rect 34296 1408 34302 1420
rect 35986 1408 35992 1420
rect 34296 1380 35992 1408
rect 34296 1368 34302 1380
rect 35986 1368 35992 1380
rect 36044 1368 36050 1420
<< via1 >>
rect 2136 48152 2188 48204
rect 14004 48152 14056 48204
rect 3608 48084 3660 48136
rect 13176 48084 13228 48136
rect 3792 48016 3844 48068
rect 15108 48016 15160 48068
rect 12992 47948 13044 48000
rect 22468 47948 22520 48000
rect 10416 47880 10468 47932
rect 20260 47880 20312 47932
rect 6368 47744 6420 47796
rect 17500 47744 17552 47796
rect 5080 47676 5132 47728
rect 16304 47676 16356 47728
rect 1400 47608 1452 47660
rect 12072 47608 12124 47660
rect 12716 47608 12768 47660
rect 27528 47608 27580 47660
rect 8944 47540 8996 47592
rect 19984 47540 20036 47592
rect 5264 47472 5316 47524
rect 17132 47472 17184 47524
rect 7104 47404 7156 47456
rect 13912 47404 13964 47456
rect 20536 47404 20588 47456
rect 30748 47404 30800 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 388 47200 440 47252
rect 2320 47200 2372 47252
rect 4620 47200 4672 47252
rect 6552 47243 6604 47252
rect 6552 47209 6561 47243
rect 6561 47209 6595 47243
rect 6595 47209 6604 47243
rect 6552 47200 6604 47209
rect 7288 47243 7340 47252
rect 7288 47209 7297 47243
rect 7297 47209 7331 47243
rect 7331 47209 7340 47243
rect 7288 47200 7340 47209
rect 8116 47243 8168 47252
rect 8116 47209 8125 47243
rect 8125 47209 8159 47243
rect 8159 47209 8168 47243
rect 8116 47200 8168 47209
rect 8668 47200 8720 47252
rect 9680 47200 9732 47252
rect 10600 47243 10652 47252
rect 10600 47209 10609 47243
rect 10609 47209 10643 47243
rect 10643 47209 10652 47243
rect 10600 47200 10652 47209
rect 11152 47200 11204 47252
rect 12440 47243 12492 47252
rect 12440 47209 12449 47243
rect 12449 47209 12483 47243
rect 12483 47209 12492 47243
rect 12440 47200 12492 47209
rect 12808 47200 12860 47252
rect 13820 47200 13872 47252
rect 14556 47200 14608 47252
rect 15384 47200 15436 47252
rect 17040 47200 17092 47252
rect 17960 47200 18012 47252
rect 19524 47200 19576 47252
rect 20720 47200 20772 47252
rect 22100 47200 22152 47252
rect 23112 47243 23164 47252
rect 23112 47209 23121 47243
rect 23121 47209 23155 47243
rect 23155 47209 23164 47243
rect 23112 47200 23164 47209
rect 23664 47200 23716 47252
rect 25320 47200 25372 47252
rect 27528 47243 27580 47252
rect 27528 47209 27537 47243
rect 27537 47209 27571 47243
rect 27571 47209 27580 47243
rect 27528 47200 27580 47209
rect 30748 47200 30800 47252
rect 3976 47132 4028 47184
rect 1400 47039 1452 47048
rect 1400 47005 1409 47039
rect 1409 47005 1443 47039
rect 1443 47005 1452 47039
rect 1400 46996 1452 47005
rect 2136 47039 2188 47048
rect 2136 47005 2145 47039
rect 2145 47005 2179 47039
rect 2179 47005 2188 47039
rect 2136 46996 2188 47005
rect 3608 46996 3660 47048
rect 3792 47039 3844 47048
rect 3792 47005 3801 47039
rect 3801 47005 3835 47039
rect 3835 47005 3844 47039
rect 3792 46996 3844 47005
rect 5080 46996 5132 47048
rect 5264 47039 5316 47048
rect 5264 47005 5273 47039
rect 5273 47005 5307 47039
rect 5307 47005 5316 47039
rect 5264 46996 5316 47005
rect 6368 47039 6420 47048
rect 6368 47005 6377 47039
rect 6377 47005 6411 47039
rect 6411 47005 6420 47039
rect 6368 46996 6420 47005
rect 7104 47039 7156 47048
rect 7104 47005 7113 47039
rect 7113 47005 7147 47039
rect 7147 47005 7156 47039
rect 7104 46996 7156 47005
rect 8944 47039 8996 47048
rect 1216 46928 1268 46980
rect 2964 46928 3016 46980
rect 8944 47005 8953 47039
rect 8953 47005 8987 47039
rect 8987 47005 8996 47039
rect 8944 46996 8996 47005
rect 21088 47132 21140 47184
rect 31024 47132 31076 47184
rect 10416 47039 10468 47048
rect 10416 47005 10425 47039
rect 10425 47005 10459 47039
rect 10459 47005 10468 47039
rect 10416 46996 10468 47005
rect 11520 47039 11572 47048
rect 11520 47005 11529 47039
rect 11529 47005 11563 47039
rect 11563 47005 11572 47039
rect 11520 46996 11572 47005
rect 12992 47039 13044 47048
rect 12992 47005 13001 47039
rect 13001 47005 13035 47039
rect 13035 47005 13044 47039
rect 12992 46996 13044 47005
rect 13268 46996 13320 47048
rect 14832 47039 14884 47048
rect 14832 47005 14841 47039
rect 14841 47005 14875 47039
rect 14875 47005 14884 47039
rect 14832 46996 14884 47005
rect 15568 47039 15620 47048
rect 15568 47005 15577 47039
rect 15577 47005 15611 47039
rect 15611 47005 15620 47039
rect 15568 46996 15620 47005
rect 16580 46996 16632 47048
rect 28172 47064 28224 47116
rect 29000 47064 29052 47116
rect 35900 47107 35952 47116
rect 35900 47073 35909 47107
rect 35909 47073 35943 47107
rect 35943 47073 35952 47107
rect 35900 47064 35952 47073
rect 37832 47064 37884 47116
rect 17408 47039 17460 47048
rect 17408 47005 17417 47039
rect 17417 47005 17451 47039
rect 17451 47005 17460 47039
rect 17408 46996 17460 47005
rect 18144 47039 18196 47048
rect 18144 47005 18153 47039
rect 18153 47005 18187 47039
rect 18187 47005 18196 47039
rect 18144 46996 18196 47005
rect 18236 46996 18288 47048
rect 19340 46996 19392 47048
rect 20720 47039 20772 47048
rect 20720 47005 20729 47039
rect 20729 47005 20763 47039
rect 20763 47005 20772 47039
rect 20720 46996 20772 47005
rect 22100 47039 22152 47048
rect 22100 47005 22109 47039
rect 22109 47005 22143 47039
rect 22143 47005 22152 47039
rect 22100 46996 22152 47005
rect 22928 47039 22980 47048
rect 22928 47005 22937 47039
rect 22937 47005 22971 47039
rect 22971 47005 22980 47039
rect 22928 46996 22980 47005
rect 24400 47039 24452 47048
rect 24400 47005 24409 47039
rect 24409 47005 24443 47039
rect 24443 47005 24452 47039
rect 24400 46996 24452 47005
rect 16212 46860 16264 46912
rect 23388 46928 23440 46980
rect 23940 46928 23992 46980
rect 24584 46928 24636 46980
rect 27068 46996 27120 47048
rect 29828 47039 29880 47048
rect 29828 47005 29837 47039
rect 29837 47005 29871 47039
rect 29871 47005 29880 47039
rect 29828 46996 29880 47005
rect 31484 47039 31536 47048
rect 31484 47005 31493 47039
rect 31493 47005 31527 47039
rect 31527 47005 31536 47039
rect 31484 46996 31536 47005
rect 27896 46928 27948 46980
rect 18052 46860 18104 46912
rect 18696 46860 18748 46912
rect 24492 46860 24544 46912
rect 30380 46860 30432 46912
rect 32404 47039 32456 47048
rect 32404 47005 32413 47039
rect 32413 47005 32447 47039
rect 32447 47005 32456 47039
rect 32404 46996 32456 47005
rect 33876 47039 33928 47048
rect 33876 47005 33885 47039
rect 33885 47005 33919 47039
rect 33919 47005 33928 47039
rect 33876 46996 33928 47005
rect 35348 46996 35400 47048
rect 36176 47039 36228 47048
rect 36176 47005 36185 47039
rect 36185 47005 36219 47039
rect 36219 47005 36228 47039
rect 36176 46996 36228 47005
rect 37556 47039 37608 47048
rect 37556 47005 37565 47039
rect 37565 47005 37599 47039
rect 37599 47005 37608 47039
rect 37556 46996 37608 47005
rect 34060 46971 34112 46980
rect 34060 46937 34069 46971
rect 34069 46937 34103 46971
rect 34103 46937 34112 46971
rect 34060 46928 34112 46937
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 5356 46656 5408 46708
rect 13268 46656 13320 46708
rect 15568 46656 15620 46708
rect 17408 46656 17460 46708
rect 18236 46656 18288 46708
rect 19340 46656 19392 46708
rect 20720 46656 20772 46708
rect 22100 46656 22152 46708
rect 5448 46563 5500 46572
rect 5448 46529 5457 46563
rect 5457 46529 5491 46563
rect 5491 46529 5500 46563
rect 5448 46520 5500 46529
rect 12256 46520 12308 46572
rect 14004 46520 14056 46572
rect 14464 46563 14516 46572
rect 14464 46529 14473 46563
rect 14473 46529 14507 46563
rect 14507 46529 14516 46563
rect 14464 46520 14516 46529
rect 16488 46520 16540 46572
rect 21364 46588 21416 46640
rect 26148 46656 26200 46708
rect 34704 46631 34756 46640
rect 11704 46452 11756 46504
rect 15108 46452 15160 46504
rect 17868 46563 17920 46572
rect 17868 46529 17877 46563
rect 17877 46529 17911 46563
rect 17911 46529 17920 46563
rect 17868 46520 17920 46529
rect 18696 46563 18748 46572
rect 18696 46529 18705 46563
rect 18705 46529 18739 46563
rect 18739 46529 18748 46563
rect 18696 46520 18748 46529
rect 17776 46452 17828 46504
rect 14832 46384 14884 46436
rect 16580 46384 16632 46436
rect 21180 46563 21232 46572
rect 21180 46529 21189 46563
rect 21189 46529 21223 46563
rect 21223 46529 21232 46563
rect 21180 46520 21232 46529
rect 24032 46563 24084 46572
rect 19340 46452 19392 46504
rect 24032 46529 24041 46563
rect 24041 46529 24075 46563
rect 24075 46529 24084 46563
rect 24032 46520 24084 46529
rect 34704 46597 34713 46631
rect 34713 46597 34747 46631
rect 34747 46597 34756 46631
rect 34704 46588 34756 46597
rect 29644 46563 29696 46572
rect 29644 46529 29653 46563
rect 29653 46529 29687 46563
rect 29687 46529 29696 46563
rect 29644 46520 29696 46529
rect 32312 46563 32364 46572
rect 32312 46529 32321 46563
rect 32321 46529 32355 46563
rect 32355 46529 32364 46563
rect 32312 46520 32364 46529
rect 32864 46520 32916 46572
rect 38660 46520 38712 46572
rect 29920 46495 29972 46504
rect 29920 46461 29929 46495
rect 29929 46461 29963 46495
rect 29963 46461 29972 46495
rect 29920 46452 29972 46461
rect 37464 46452 37516 46504
rect 14924 46316 14976 46368
rect 21272 46384 21324 46436
rect 32128 46359 32180 46368
rect 32128 46325 32137 46359
rect 32137 46325 32171 46359
rect 32171 46325 32180 46359
rect 32128 46316 32180 46325
rect 32956 46359 33008 46368
rect 32956 46325 32965 46359
rect 32965 46325 32999 46359
rect 32999 46325 33008 46359
rect 32956 46316 33008 46325
rect 34796 46359 34848 46368
rect 34796 46325 34805 46359
rect 34805 46325 34839 46359
rect 34839 46325 34848 46359
rect 34796 46316 34848 46325
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 5448 46112 5500 46164
rect 12256 46155 12308 46164
rect 12256 46121 12265 46155
rect 12265 46121 12299 46155
rect 12299 46121 12308 46155
rect 12256 46112 12308 46121
rect 14464 46112 14516 46164
rect 14924 46112 14976 46164
rect 16488 46155 16540 46164
rect 16488 46121 16497 46155
rect 16497 46121 16531 46155
rect 16531 46121 16540 46155
rect 16488 46112 16540 46121
rect 18144 46112 18196 46164
rect 22928 46112 22980 46164
rect 17868 46044 17920 46096
rect 10692 45976 10744 46028
rect 14096 45976 14148 46028
rect 11980 45951 12032 45960
rect 11980 45917 11989 45951
rect 11989 45917 12023 45951
rect 12023 45917 12032 45951
rect 11980 45908 12032 45917
rect 12072 45951 12124 45960
rect 12072 45917 12081 45951
rect 12081 45917 12115 45951
rect 12115 45917 12124 45951
rect 13268 45951 13320 45960
rect 12072 45908 12124 45917
rect 13268 45917 13277 45951
rect 13277 45917 13311 45951
rect 13311 45917 13320 45951
rect 13268 45908 13320 45917
rect 14464 45951 14516 45960
rect 14464 45917 14473 45951
rect 14473 45917 14507 45951
rect 14507 45917 14516 45951
rect 14464 45908 14516 45917
rect 15108 45976 15160 46028
rect 15476 45951 15528 45960
rect 13912 45840 13964 45892
rect 15476 45917 15485 45951
rect 15485 45917 15519 45951
rect 15519 45917 15528 45951
rect 15476 45908 15528 45917
rect 16304 45951 16356 45960
rect 16304 45917 16313 45951
rect 16313 45917 16347 45951
rect 16347 45917 16356 45951
rect 23296 45976 23348 46028
rect 16304 45908 16356 45917
rect 17132 45951 17184 45960
rect 17132 45917 17141 45951
rect 17141 45917 17175 45951
rect 17175 45917 17184 45951
rect 17132 45908 17184 45917
rect 22376 45951 22428 45960
rect 22376 45917 22385 45951
rect 22385 45917 22419 45951
rect 22419 45917 22428 45951
rect 22376 45908 22428 45917
rect 37188 45951 37240 45960
rect 37188 45917 37197 45951
rect 37197 45917 37231 45951
rect 37231 45917 37240 45951
rect 37188 45908 37240 45917
rect 39488 45908 39540 45960
rect 17224 45840 17276 45892
rect 15476 45772 15528 45824
rect 37280 45815 37332 45824
rect 37280 45781 37289 45815
rect 37289 45781 37323 45815
rect 37323 45781 37332 45815
rect 37280 45772 37332 45781
rect 38016 45815 38068 45824
rect 38016 45781 38025 45815
rect 38025 45781 38059 45815
rect 38059 45781 38068 45815
rect 38016 45772 38068 45781
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 13268 45568 13320 45620
rect 18144 45568 18196 45620
rect 23296 45611 23348 45620
rect 23296 45577 23305 45611
rect 23305 45577 23339 45611
rect 23339 45577 23348 45611
rect 23296 45568 23348 45577
rect 18696 45500 18748 45552
rect 21180 45500 21232 45552
rect 22376 45500 22428 45552
rect 24032 45500 24084 45552
rect 12256 45432 12308 45484
rect 14004 45432 14056 45484
rect 17500 45475 17552 45484
rect 17500 45441 17509 45475
rect 17509 45441 17543 45475
rect 17543 45441 17552 45475
rect 17500 45432 17552 45441
rect 18328 45432 18380 45484
rect 19984 45475 20036 45484
rect 19984 45441 19993 45475
rect 19993 45441 20027 45475
rect 20027 45441 20036 45475
rect 19984 45432 20036 45441
rect 21088 45475 21140 45484
rect 21088 45441 21097 45475
rect 21097 45441 21131 45475
rect 21131 45441 21140 45475
rect 21088 45432 21140 45441
rect 22468 45475 22520 45484
rect 22468 45441 22477 45475
rect 22477 45441 22511 45475
rect 22511 45441 22520 45475
rect 22468 45432 22520 45441
rect 24216 45432 24268 45484
rect 30380 45432 30432 45484
rect 13544 45407 13596 45416
rect 13544 45373 13553 45407
rect 13553 45373 13587 45407
rect 13587 45373 13596 45407
rect 13544 45364 13596 45373
rect 17316 45407 17368 45416
rect 17316 45373 17325 45407
rect 17325 45373 17359 45407
rect 17359 45373 17368 45407
rect 17316 45364 17368 45373
rect 20628 45364 20680 45416
rect 22928 45364 22980 45416
rect 13912 45296 13964 45348
rect 19340 45296 19392 45348
rect 21088 45296 21140 45348
rect 15476 45228 15528 45280
rect 22928 45271 22980 45280
rect 22928 45237 22937 45271
rect 22937 45237 22971 45271
rect 22971 45237 22980 45271
rect 22928 45228 22980 45237
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 21364 45067 21416 45076
rect 21364 45033 21373 45067
rect 21373 45033 21407 45067
rect 21407 45033 21416 45067
rect 21364 45024 21416 45033
rect 17500 44956 17552 45008
rect 25044 44956 25096 45008
rect 18696 44888 18748 44940
rect 19984 44888 20036 44940
rect 22468 44888 22520 44940
rect 18144 44863 18196 44872
rect 18144 44829 18153 44863
rect 18153 44829 18187 44863
rect 18187 44829 18196 44863
rect 18144 44820 18196 44829
rect 19248 44820 19300 44872
rect 23020 44863 23072 44872
rect 23020 44829 23029 44863
rect 23029 44829 23063 44863
rect 23063 44829 23072 44863
rect 23020 44820 23072 44829
rect 21732 44752 21784 44804
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 16856 44480 16908 44532
rect 17316 44480 17368 44532
rect 18328 44523 18380 44532
rect 18328 44489 18337 44523
rect 18337 44489 18371 44523
rect 18371 44489 18380 44523
rect 18328 44480 18380 44489
rect 24400 44480 24452 44532
rect 14556 44344 14608 44396
rect 14832 44344 14884 44396
rect 18052 44344 18104 44396
rect 20076 44387 20128 44396
rect 20076 44353 20110 44387
rect 20110 44353 20128 44387
rect 20076 44344 20128 44353
rect 20996 44344 21048 44396
rect 24032 44387 24084 44396
rect 24032 44353 24041 44387
rect 24041 44353 24075 44387
rect 24075 44353 24084 44387
rect 24032 44344 24084 44353
rect 12900 44319 12952 44328
rect 12900 44285 12909 44319
rect 12909 44285 12943 44319
rect 12943 44285 12952 44319
rect 12900 44276 12952 44285
rect 14648 44276 14700 44328
rect 19800 44319 19852 44328
rect 19800 44285 19809 44319
rect 19809 44285 19843 44319
rect 19843 44285 19852 44319
rect 19800 44276 19852 44285
rect 23480 44276 23532 44328
rect 18144 44208 18196 44260
rect 14464 44140 14516 44192
rect 21088 44140 21140 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 19984 43936 20036 43988
rect 20628 43979 20680 43988
rect 20628 43945 20637 43979
rect 20637 43945 20671 43979
rect 20671 43945 20680 43979
rect 20628 43936 20680 43945
rect 20260 43868 20312 43920
rect 22652 43936 22704 43988
rect 24032 43936 24084 43988
rect 18052 43800 18104 43852
rect 14464 43732 14516 43784
rect 14648 43732 14700 43784
rect 16672 43732 16724 43784
rect 17500 43775 17552 43784
rect 17500 43741 17509 43775
rect 17509 43741 17543 43775
rect 17543 43741 17552 43775
rect 17500 43732 17552 43741
rect 19800 43732 19852 43784
rect 22008 43732 22060 43784
rect 15016 43596 15068 43648
rect 15292 43664 15344 43716
rect 19340 43664 19392 43716
rect 20720 43664 20772 43716
rect 15384 43596 15436 43648
rect 17224 43596 17276 43648
rect 22100 43596 22152 43648
rect 22652 43707 22704 43716
rect 22652 43673 22661 43707
rect 22661 43673 22695 43707
rect 22695 43673 22704 43707
rect 23296 43732 23348 43784
rect 22652 43664 22704 43673
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 14096 43435 14148 43444
rect 14096 43401 14105 43435
rect 14105 43401 14139 43435
rect 14139 43401 14148 43435
rect 14096 43392 14148 43401
rect 14556 43435 14608 43444
rect 14556 43401 14565 43435
rect 14565 43401 14599 43435
rect 14599 43401 14608 43435
rect 14556 43392 14608 43401
rect 23940 43435 23992 43444
rect 23940 43401 23949 43435
rect 23949 43401 23983 43435
rect 23983 43401 23992 43435
rect 23940 43392 23992 43401
rect 24584 43435 24636 43444
rect 24584 43401 24593 43435
rect 24593 43401 24627 43435
rect 24627 43401 24636 43435
rect 24584 43392 24636 43401
rect 14648 43324 14700 43376
rect 21088 43324 21140 43376
rect 14096 43256 14148 43308
rect 14924 43299 14976 43308
rect 14924 43265 14933 43299
rect 14933 43265 14967 43299
rect 14967 43265 14976 43299
rect 14924 43256 14976 43265
rect 15016 43299 15068 43308
rect 15016 43265 15025 43299
rect 15025 43265 15059 43299
rect 15059 43265 15068 43299
rect 15200 43299 15252 43308
rect 15016 43256 15068 43265
rect 15200 43265 15209 43299
rect 15209 43265 15243 43299
rect 15243 43265 15252 43299
rect 15200 43256 15252 43265
rect 15384 43256 15436 43308
rect 16672 43299 16724 43308
rect 15936 43120 15988 43172
rect 16028 43052 16080 43104
rect 16672 43265 16681 43299
rect 16681 43265 16715 43299
rect 16715 43265 16724 43299
rect 16672 43256 16724 43265
rect 16764 43256 16816 43308
rect 19892 43299 19944 43308
rect 19892 43265 19901 43299
rect 19901 43265 19935 43299
rect 19935 43265 19944 43299
rect 19892 43256 19944 43265
rect 24124 43299 24176 43308
rect 24124 43265 24133 43299
rect 24133 43265 24167 43299
rect 24167 43265 24176 43299
rect 24124 43256 24176 43265
rect 24768 43299 24820 43308
rect 24768 43265 24777 43299
rect 24777 43265 24811 43299
rect 24811 43265 24820 43299
rect 24768 43256 24820 43265
rect 18144 43052 18196 43104
rect 20628 43052 20680 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 16764 42848 16816 42900
rect 24768 42891 24820 42900
rect 24768 42857 24777 42891
rect 24777 42857 24811 42891
rect 24811 42857 24820 42891
rect 24768 42848 24820 42857
rect 20720 42780 20772 42832
rect 20904 42780 20956 42832
rect 14096 42755 14148 42764
rect 14096 42721 14105 42755
rect 14105 42721 14139 42755
rect 14139 42721 14148 42755
rect 14096 42712 14148 42721
rect 14188 42712 14240 42764
rect 14004 42644 14056 42696
rect 14372 42687 14424 42696
rect 14372 42653 14381 42687
rect 14381 42653 14415 42687
rect 14415 42653 14424 42687
rect 14372 42644 14424 42653
rect 14924 42712 14976 42764
rect 14740 42687 14792 42696
rect 13268 42576 13320 42628
rect 14740 42653 14749 42687
rect 14749 42653 14783 42687
rect 14783 42653 14792 42687
rect 14740 42644 14792 42653
rect 15200 42644 15252 42696
rect 16028 42687 16080 42696
rect 16028 42653 16037 42687
rect 16037 42653 16071 42687
rect 16071 42653 16080 42687
rect 16028 42644 16080 42653
rect 16212 42687 16264 42696
rect 16212 42653 16221 42687
rect 16221 42653 16255 42687
rect 16255 42653 16264 42687
rect 16212 42644 16264 42653
rect 19984 42644 20036 42696
rect 20260 42644 20312 42696
rect 23388 42712 23440 42764
rect 21180 42687 21232 42696
rect 17408 42576 17460 42628
rect 19892 42576 19944 42628
rect 14004 42508 14056 42560
rect 14924 42508 14976 42560
rect 19432 42508 19484 42560
rect 20720 42576 20772 42628
rect 21180 42653 21189 42687
rect 21189 42653 21223 42687
rect 21223 42653 21232 42687
rect 21180 42644 21232 42653
rect 27712 42712 27764 42764
rect 20444 42508 20496 42560
rect 22100 42576 22152 42628
rect 22652 42619 22704 42628
rect 22652 42585 22661 42619
rect 22661 42585 22695 42619
rect 22695 42585 22704 42619
rect 22652 42576 22704 42585
rect 22836 42551 22888 42560
rect 22836 42517 22845 42551
rect 22845 42517 22879 42551
rect 22879 42517 22888 42551
rect 22836 42508 22888 42517
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 14832 42304 14884 42356
rect 15292 42347 15344 42356
rect 15292 42313 15301 42347
rect 15301 42313 15335 42347
rect 15335 42313 15344 42347
rect 15292 42304 15344 42313
rect 17500 42347 17552 42356
rect 17500 42313 17509 42347
rect 17509 42313 17543 42347
rect 17543 42313 17552 42347
rect 17500 42304 17552 42313
rect 19340 42304 19392 42356
rect 20076 42304 20128 42356
rect 24124 42304 24176 42356
rect 14280 42168 14332 42220
rect 16304 42236 16356 42288
rect 14832 42211 14884 42220
rect 14188 42100 14240 42152
rect 14832 42177 14841 42211
rect 14841 42177 14875 42211
rect 14875 42177 14884 42211
rect 14832 42168 14884 42177
rect 15568 42168 15620 42220
rect 15844 42168 15896 42220
rect 14372 41964 14424 42016
rect 14740 41964 14792 42016
rect 14832 41964 14884 42016
rect 16120 42168 16172 42220
rect 18052 42168 18104 42220
rect 16212 42100 16264 42152
rect 17316 42075 17368 42084
rect 17316 42041 17325 42075
rect 17325 42041 17359 42075
rect 17359 42041 17368 42075
rect 17316 42032 17368 42041
rect 19524 42211 19576 42220
rect 19524 42177 19533 42211
rect 19533 42177 19567 42211
rect 19567 42177 19576 42211
rect 19524 42168 19576 42177
rect 20352 42168 20404 42220
rect 20904 42236 20956 42288
rect 20628 42211 20680 42220
rect 20628 42177 20637 42211
rect 20637 42177 20671 42211
rect 20671 42177 20680 42211
rect 20628 42168 20680 42177
rect 20812 42211 20864 42220
rect 20812 42177 20821 42211
rect 20821 42177 20855 42211
rect 20855 42177 20864 42211
rect 20812 42168 20864 42177
rect 21180 42168 21232 42220
rect 22008 42211 22060 42220
rect 22008 42177 22017 42211
rect 22017 42177 22051 42211
rect 22051 42177 22060 42211
rect 22008 42168 22060 42177
rect 21456 42100 21508 42152
rect 24032 42211 24084 42220
rect 24032 42177 24041 42211
rect 24041 42177 24075 42211
rect 24075 42177 24084 42211
rect 24032 42168 24084 42177
rect 27528 42168 27580 42220
rect 23848 42143 23900 42152
rect 23848 42109 23857 42143
rect 23857 42109 23891 42143
rect 23891 42109 23900 42143
rect 23848 42100 23900 42109
rect 19984 42032 20036 42084
rect 17960 42007 18012 42016
rect 17960 41973 17969 42007
rect 17969 41973 18003 42007
rect 18003 41973 18012 42007
rect 17960 41964 18012 41973
rect 20260 41964 20312 42016
rect 20444 41964 20496 42016
rect 22652 41964 22704 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 11520 41760 11572 41812
rect 16672 41760 16724 41812
rect 17684 41760 17736 41812
rect 22008 41760 22060 41812
rect 27528 41803 27580 41812
rect 27528 41769 27537 41803
rect 27537 41769 27571 41803
rect 27571 41769 27580 41803
rect 27528 41760 27580 41769
rect 24032 41692 24084 41744
rect 14188 41624 14240 41676
rect 15292 41624 15344 41676
rect 15844 41624 15896 41676
rect 13268 41420 13320 41472
rect 13452 41420 13504 41472
rect 20904 41556 20956 41608
rect 21180 41556 21232 41608
rect 14556 41488 14608 41540
rect 15200 41488 15252 41540
rect 27252 41488 27304 41540
rect 27988 41488 28040 41540
rect 19340 41420 19392 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 13268 41216 13320 41268
rect 13176 41148 13228 41200
rect 15292 41216 15344 41268
rect 15568 41216 15620 41268
rect 15384 41148 15436 41200
rect 16856 41216 16908 41268
rect 18052 41216 18104 41268
rect 18328 41216 18380 41268
rect 34060 41216 34112 41268
rect 13268 41080 13320 41132
rect 15844 41148 15896 41200
rect 16212 41148 16264 41200
rect 17040 41191 17092 41200
rect 17040 41157 17049 41191
rect 17049 41157 17083 41191
rect 17083 41157 17092 41191
rect 17040 41148 17092 41157
rect 17960 41191 18012 41200
rect 17960 41157 17994 41191
rect 17994 41157 18012 41191
rect 17960 41148 18012 41157
rect 18236 41148 18288 41200
rect 21640 41148 21692 41200
rect 21824 41148 21876 41200
rect 22284 41148 22336 41200
rect 34796 41148 34848 41200
rect 17684 41123 17736 41132
rect 12992 41012 13044 41064
rect 13728 41012 13780 41064
rect 14832 41012 14884 41064
rect 17684 41089 17693 41123
rect 17693 41089 17727 41123
rect 17727 41089 17736 41123
rect 17684 41080 17736 41089
rect 18328 41080 18380 41132
rect 22008 41080 22060 41132
rect 19524 41055 19576 41064
rect 19524 41021 19533 41055
rect 19533 41021 19567 41055
rect 19567 41021 19576 41055
rect 19524 41012 19576 41021
rect 13452 40944 13504 40996
rect 17316 40944 17368 40996
rect 17592 40944 17644 40996
rect 20812 41012 20864 41064
rect 21364 41012 21416 41064
rect 21916 41055 21968 41064
rect 21916 41021 21925 41055
rect 21925 41021 21959 41055
rect 21959 41021 21968 41055
rect 21916 41012 21968 41021
rect 20444 40944 20496 40996
rect 13084 40919 13136 40928
rect 13084 40885 13093 40919
rect 13093 40885 13127 40919
rect 13127 40885 13136 40919
rect 13084 40876 13136 40885
rect 13268 40876 13320 40928
rect 15844 40876 15896 40928
rect 15936 40919 15988 40928
rect 15936 40885 15945 40919
rect 15945 40885 15979 40919
rect 15979 40885 15988 40919
rect 15936 40876 15988 40885
rect 18328 40876 18380 40928
rect 21548 40876 21600 40928
rect 23848 40944 23900 40996
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 12256 40715 12308 40724
rect 12256 40681 12265 40715
rect 12265 40681 12299 40715
rect 12299 40681 12308 40715
rect 12256 40672 12308 40681
rect 13084 40715 13136 40724
rect 13084 40681 13093 40715
rect 13093 40681 13127 40715
rect 13127 40681 13136 40715
rect 13084 40672 13136 40681
rect 16304 40672 16356 40724
rect 17040 40672 17092 40724
rect 21456 40672 21508 40724
rect 21640 40672 21692 40724
rect 25412 40672 25464 40724
rect 16396 40604 16448 40656
rect 19524 40604 19576 40656
rect 14648 40579 14700 40588
rect 14648 40545 14657 40579
rect 14657 40545 14691 40579
rect 14691 40545 14700 40579
rect 14648 40536 14700 40545
rect 12532 40468 12584 40520
rect 15936 40468 15988 40520
rect 13176 40400 13228 40452
rect 14924 40443 14976 40452
rect 14924 40409 14958 40443
rect 14958 40409 14976 40443
rect 14924 40400 14976 40409
rect 13084 40375 13136 40384
rect 13084 40341 13093 40375
rect 13093 40341 13127 40375
rect 13127 40341 13136 40375
rect 13084 40332 13136 40341
rect 13268 40375 13320 40384
rect 13268 40341 13277 40375
rect 13277 40341 13311 40375
rect 13311 40341 13320 40375
rect 13268 40332 13320 40341
rect 16948 40536 17000 40588
rect 16488 40511 16540 40520
rect 16488 40477 16497 40511
rect 16497 40477 16531 40511
rect 16531 40477 16540 40511
rect 16488 40468 16540 40477
rect 16764 40468 16816 40520
rect 17316 40511 17368 40520
rect 17316 40477 17325 40511
rect 17325 40477 17359 40511
rect 17359 40477 17368 40511
rect 17316 40468 17368 40477
rect 17960 40511 18012 40520
rect 17960 40477 17969 40511
rect 17969 40477 18003 40511
rect 18003 40477 18012 40511
rect 17960 40468 18012 40477
rect 19340 40468 19392 40520
rect 20812 40468 20864 40520
rect 21180 40536 21232 40588
rect 21364 40468 21416 40520
rect 17592 40400 17644 40452
rect 21824 40443 21876 40452
rect 16580 40332 16632 40384
rect 16856 40332 16908 40384
rect 17224 40332 17276 40384
rect 18788 40332 18840 40384
rect 20260 40332 20312 40384
rect 21824 40409 21833 40443
rect 21833 40409 21867 40443
rect 21867 40409 21876 40443
rect 21824 40400 21876 40409
rect 22008 40468 22060 40520
rect 22284 40511 22336 40520
rect 22284 40477 22298 40511
rect 22298 40477 22332 40511
rect 22332 40477 22336 40511
rect 22284 40468 22336 40477
rect 22836 40332 22888 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 13268 40060 13320 40112
rect 17868 40128 17920 40180
rect 19248 40171 19300 40180
rect 19248 40137 19257 40171
rect 19257 40137 19291 40171
rect 19291 40137 19300 40171
rect 19248 40128 19300 40137
rect 12072 39992 12124 40044
rect 12900 39992 12952 40044
rect 16948 40060 17000 40112
rect 11520 39967 11572 39976
rect 11520 39933 11529 39967
rect 11529 39933 11563 39967
rect 11563 39933 11572 39967
rect 11520 39924 11572 39933
rect 17224 39992 17276 40044
rect 18512 40035 18564 40044
rect 18512 40001 18521 40035
rect 18521 40001 18555 40035
rect 18555 40001 18564 40035
rect 18512 39992 18564 40001
rect 20260 40060 20312 40112
rect 21548 40060 21600 40112
rect 23204 40128 23256 40180
rect 25504 40060 25556 40112
rect 15108 39924 15160 39976
rect 17316 39924 17368 39976
rect 17960 39924 18012 39976
rect 22284 39992 22336 40044
rect 24860 40035 24912 40044
rect 24860 40001 24869 40035
rect 24869 40001 24903 40035
rect 24903 40001 24912 40035
rect 24860 39992 24912 40001
rect 25044 40035 25096 40044
rect 25044 40001 25053 40035
rect 25053 40001 25087 40035
rect 25087 40001 25096 40035
rect 25044 39992 25096 40001
rect 23204 39924 23256 39976
rect 15660 39856 15712 39908
rect 16304 39856 16356 39908
rect 19340 39856 19392 39908
rect 14188 39831 14240 39840
rect 14188 39797 14197 39831
rect 14197 39797 14231 39831
rect 14231 39797 14240 39831
rect 14188 39788 14240 39797
rect 15384 39788 15436 39840
rect 20536 39856 20588 39908
rect 23296 39899 23348 39908
rect 23296 39865 23305 39899
rect 23305 39865 23339 39899
rect 23339 39865 23348 39899
rect 23296 39856 23348 39865
rect 23480 39899 23532 39908
rect 23480 39865 23489 39899
rect 23489 39865 23523 39899
rect 23523 39865 23532 39899
rect 23480 39856 23532 39865
rect 20260 39831 20312 39840
rect 20260 39797 20269 39831
rect 20269 39797 20303 39831
rect 20303 39797 20312 39831
rect 20260 39788 20312 39797
rect 24308 39831 24360 39840
rect 24308 39797 24317 39831
rect 24317 39797 24351 39831
rect 24351 39797 24360 39831
rect 24308 39788 24360 39797
rect 36176 39788 36228 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 12532 39627 12584 39636
rect 12532 39593 12541 39627
rect 12541 39593 12575 39627
rect 12575 39593 12584 39627
rect 12532 39584 12584 39593
rect 13084 39584 13136 39636
rect 14924 39627 14976 39636
rect 14924 39593 14933 39627
rect 14933 39593 14967 39627
rect 14967 39593 14976 39627
rect 14924 39584 14976 39593
rect 12256 39380 12308 39432
rect 12624 39380 12676 39432
rect 16764 39584 16816 39636
rect 24860 39584 24912 39636
rect 25412 39584 25464 39636
rect 25136 39559 25188 39568
rect 25136 39525 25145 39559
rect 25145 39525 25179 39559
rect 25179 39525 25188 39559
rect 25136 39516 25188 39525
rect 15660 39448 15712 39500
rect 15936 39448 15988 39500
rect 14280 39312 14332 39364
rect 15384 39423 15436 39432
rect 15384 39389 15393 39423
rect 15393 39389 15427 39423
rect 15427 39389 15436 39423
rect 15384 39380 15436 39389
rect 15844 39380 15896 39432
rect 19432 39423 19484 39432
rect 19432 39389 19441 39423
rect 19441 39389 19475 39423
rect 19475 39389 19484 39423
rect 19432 39380 19484 39389
rect 21088 39380 21140 39432
rect 21916 39423 21968 39432
rect 21916 39389 21925 39423
rect 21925 39389 21959 39423
rect 21959 39389 21968 39423
rect 21916 39380 21968 39389
rect 32956 39584 33008 39636
rect 15476 39312 15528 39364
rect 17868 39355 17920 39364
rect 17868 39321 17877 39355
rect 17877 39321 17911 39355
rect 17911 39321 17920 39355
rect 17868 39312 17920 39321
rect 18512 39312 18564 39364
rect 20996 39355 21048 39364
rect 20996 39321 21005 39355
rect 21005 39321 21039 39355
rect 21039 39321 21048 39355
rect 20996 39312 21048 39321
rect 22192 39355 22244 39364
rect 22192 39321 22226 39355
rect 22226 39321 22244 39355
rect 22192 39312 22244 39321
rect 24860 39312 24912 39364
rect 11612 39244 11664 39296
rect 15292 39244 15344 39296
rect 17224 39244 17276 39296
rect 18236 39287 18288 39296
rect 18236 39253 18245 39287
rect 18245 39253 18279 39287
rect 18279 39253 18288 39287
rect 18236 39244 18288 39253
rect 20076 39244 20128 39296
rect 20536 39287 20588 39296
rect 20536 39253 20545 39287
rect 20545 39253 20579 39287
rect 20579 39253 20588 39287
rect 20536 39244 20588 39253
rect 21456 39244 21508 39296
rect 22100 39244 22152 39296
rect 25964 39312 26016 39364
rect 26240 39287 26292 39296
rect 26240 39253 26249 39287
rect 26249 39253 26283 39287
rect 26283 39253 26292 39287
rect 26240 39244 26292 39253
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 11520 39040 11572 39092
rect 15476 39083 15528 39092
rect 15476 39049 15485 39083
rect 15485 39049 15519 39083
rect 15519 39049 15528 39083
rect 15476 39040 15528 39049
rect 15936 39040 15988 39092
rect 15660 38972 15712 39024
rect 17316 38972 17368 39024
rect 12532 38836 12584 38888
rect 15936 38947 15988 38956
rect 15936 38913 15945 38947
rect 15945 38913 15979 38947
rect 15979 38913 15988 38947
rect 21088 39040 21140 39092
rect 15936 38904 15988 38913
rect 16028 38836 16080 38888
rect 16396 38836 16448 38888
rect 11888 38811 11940 38820
rect 11888 38777 11897 38811
rect 11897 38777 11931 38811
rect 11931 38777 11940 38811
rect 11888 38768 11940 38777
rect 17592 38904 17644 38956
rect 21916 38972 21968 39024
rect 20076 38947 20128 38956
rect 20076 38913 20110 38947
rect 20110 38913 20128 38947
rect 20076 38904 20128 38913
rect 22284 38972 22336 39024
rect 26424 38947 26476 38956
rect 26424 38913 26433 38947
rect 26433 38913 26467 38947
rect 26467 38913 26476 38947
rect 26424 38904 26476 38913
rect 17684 38700 17736 38752
rect 18512 38700 18564 38752
rect 23756 38743 23808 38752
rect 23756 38709 23765 38743
rect 23765 38709 23799 38743
rect 23799 38709 23808 38743
rect 23756 38700 23808 38709
rect 25044 38700 25096 38752
rect 25320 38700 25372 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 12716 38539 12768 38548
rect 12716 38505 12725 38539
rect 12725 38505 12759 38539
rect 12759 38505 12768 38539
rect 12716 38496 12768 38505
rect 15936 38496 15988 38548
rect 17224 38496 17276 38548
rect 17592 38496 17644 38548
rect 17684 38496 17736 38548
rect 18052 38496 18104 38548
rect 20260 38496 20312 38548
rect 20812 38496 20864 38548
rect 21180 38496 21232 38548
rect 22284 38496 22336 38548
rect 23204 38539 23256 38548
rect 23204 38505 23213 38539
rect 23213 38505 23247 38539
rect 23247 38505 23256 38539
rect 23204 38496 23256 38505
rect 26240 38496 26292 38548
rect 12440 38360 12492 38412
rect 12900 38360 12952 38412
rect 15200 38360 15252 38412
rect 14280 38335 14332 38344
rect 14280 38301 14289 38335
rect 14289 38301 14323 38335
rect 14323 38301 14332 38335
rect 14280 38292 14332 38301
rect 14924 38292 14976 38344
rect 16856 38360 16908 38412
rect 17316 38360 17368 38412
rect 16948 38292 17000 38344
rect 17040 38292 17092 38344
rect 17408 38292 17460 38344
rect 18236 38360 18288 38412
rect 19432 38428 19484 38480
rect 22192 38428 22244 38480
rect 22008 38360 22060 38412
rect 12716 38224 12768 38276
rect 14648 38224 14700 38276
rect 16488 38267 16540 38276
rect 11796 38156 11848 38208
rect 12532 38156 12584 38208
rect 13452 38199 13504 38208
rect 13452 38165 13461 38199
rect 13461 38165 13495 38199
rect 13495 38165 13504 38199
rect 13452 38156 13504 38165
rect 14372 38156 14424 38208
rect 16488 38233 16497 38267
rect 16497 38233 16531 38267
rect 16531 38233 16540 38267
rect 16488 38224 16540 38233
rect 16764 38224 16816 38276
rect 16856 38199 16908 38208
rect 16856 38165 16865 38199
rect 16865 38165 16899 38199
rect 16899 38165 16908 38199
rect 16856 38156 16908 38165
rect 18052 38292 18104 38344
rect 18880 38292 18932 38344
rect 19340 38292 19392 38344
rect 17868 38224 17920 38276
rect 20076 38224 20128 38276
rect 20720 38292 20772 38344
rect 21272 38335 21324 38344
rect 21272 38301 21281 38335
rect 21281 38301 21315 38335
rect 21315 38301 21324 38335
rect 21272 38292 21324 38301
rect 20996 38224 21048 38276
rect 21456 38335 21508 38344
rect 21456 38301 21465 38335
rect 21465 38301 21499 38335
rect 21499 38301 21508 38335
rect 21456 38292 21508 38301
rect 21824 38292 21876 38344
rect 21916 38292 21968 38344
rect 22468 38428 22520 38480
rect 25136 38471 25188 38480
rect 25136 38437 25145 38471
rect 25145 38437 25179 38471
rect 25179 38437 25188 38471
rect 25136 38428 25188 38437
rect 26424 38428 26476 38480
rect 22560 38335 22612 38344
rect 22560 38301 22569 38335
rect 22569 38301 22603 38335
rect 22603 38301 22612 38335
rect 22560 38292 22612 38301
rect 23112 38292 23164 38344
rect 22836 38224 22888 38276
rect 21088 38156 21140 38208
rect 22008 38156 22060 38208
rect 23756 38292 23808 38344
rect 26056 38292 26108 38344
rect 26332 38335 26384 38344
rect 26332 38301 26341 38335
rect 26341 38301 26375 38335
rect 26375 38301 26384 38335
rect 26332 38292 26384 38301
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 10692 37995 10744 38004
rect 10692 37961 10701 37995
rect 10701 37961 10735 37995
rect 10735 37961 10744 37995
rect 10692 37952 10744 37961
rect 12348 37952 12400 38004
rect 14280 37995 14332 38004
rect 14280 37961 14289 37995
rect 14289 37961 14323 37995
rect 14323 37961 14332 37995
rect 14280 37952 14332 37961
rect 16212 37952 16264 38004
rect 16488 37952 16540 38004
rect 18420 37952 18472 38004
rect 19340 37952 19392 38004
rect 20076 37995 20128 38004
rect 20076 37961 20085 37995
rect 20085 37961 20119 37995
rect 20119 37961 20128 37995
rect 20076 37952 20128 37961
rect 21088 37952 21140 38004
rect 22560 37952 22612 38004
rect 25136 37952 25188 38004
rect 27712 37995 27764 38004
rect 27712 37961 27721 37995
rect 27721 37961 27755 37995
rect 27755 37961 27764 37995
rect 27712 37952 27764 37961
rect 28356 37952 28408 38004
rect 8944 37816 8996 37868
rect 9588 37859 9640 37868
rect 9588 37825 9622 37859
rect 9622 37825 9640 37859
rect 12440 37884 12492 37936
rect 14096 37927 14148 37936
rect 14096 37893 14105 37927
rect 14105 37893 14139 37927
rect 14139 37893 14148 37927
rect 14096 37884 14148 37893
rect 14648 37884 14700 37936
rect 9588 37816 9640 37825
rect 11612 37816 11664 37868
rect 13636 37816 13688 37868
rect 18512 37927 18564 37936
rect 18512 37893 18521 37927
rect 18521 37893 18555 37927
rect 18555 37893 18564 37927
rect 18512 37884 18564 37893
rect 16764 37748 16816 37800
rect 17868 37748 17920 37800
rect 18328 37816 18380 37868
rect 18420 37859 18472 37868
rect 18420 37825 18429 37859
rect 18429 37825 18463 37859
rect 18463 37825 18472 37859
rect 18420 37816 18472 37825
rect 18604 37859 18656 37868
rect 18604 37825 18613 37859
rect 18613 37825 18647 37859
rect 18647 37825 18656 37859
rect 20996 37884 21048 37936
rect 22100 37884 22152 37936
rect 22836 37884 22888 37936
rect 27896 37884 27948 37936
rect 18604 37816 18656 37825
rect 18512 37748 18564 37800
rect 19432 37748 19484 37800
rect 20628 37816 20680 37868
rect 20812 37816 20864 37868
rect 22008 37859 22060 37868
rect 22008 37825 22017 37859
rect 22017 37825 22051 37859
rect 22051 37825 22060 37859
rect 22008 37816 22060 37825
rect 25228 37816 25280 37868
rect 26332 37816 26384 37868
rect 26056 37748 26108 37800
rect 28356 37748 28408 37800
rect 13728 37723 13780 37732
rect 13728 37689 13737 37723
rect 13737 37689 13771 37723
rect 13771 37689 13780 37723
rect 13728 37680 13780 37689
rect 28172 37680 28224 37732
rect 28540 37723 28592 37732
rect 28540 37689 28549 37723
rect 28549 37689 28583 37723
rect 28583 37689 28592 37723
rect 28540 37680 28592 37689
rect 18236 37612 18288 37664
rect 18880 37612 18932 37664
rect 21824 37612 21876 37664
rect 37464 37680 37516 37732
rect 29552 37655 29604 37664
rect 29552 37621 29561 37655
rect 29561 37621 29595 37655
rect 29595 37621 29604 37655
rect 29552 37612 29604 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 13452 37408 13504 37460
rect 11888 37340 11940 37392
rect 13728 37340 13780 37392
rect 15660 37340 15712 37392
rect 8944 37315 8996 37324
rect 8944 37281 8953 37315
rect 8953 37281 8987 37315
rect 8987 37281 8996 37315
rect 8944 37272 8996 37281
rect 16028 37315 16080 37324
rect 16028 37281 16037 37315
rect 16037 37281 16071 37315
rect 16071 37281 16080 37315
rect 16028 37272 16080 37281
rect 13268 37204 13320 37256
rect 15752 37204 15804 37256
rect 16580 37340 16632 37392
rect 16948 37408 17000 37460
rect 18604 37408 18656 37460
rect 24308 37408 24360 37460
rect 23296 37383 23348 37392
rect 23296 37349 23305 37383
rect 23305 37349 23339 37383
rect 23339 37349 23348 37383
rect 23296 37340 23348 37349
rect 23388 37340 23440 37392
rect 17684 37315 17736 37324
rect 9404 37136 9456 37188
rect 13636 37136 13688 37188
rect 14372 37179 14424 37188
rect 14372 37145 14406 37179
rect 14406 37145 14424 37179
rect 14372 37136 14424 37145
rect 14648 37136 14700 37188
rect 16856 37204 16908 37256
rect 17684 37281 17693 37315
rect 17693 37281 17727 37315
rect 17727 37281 17736 37315
rect 17684 37272 17736 37281
rect 28908 37315 28960 37324
rect 10324 37111 10376 37120
rect 10324 37077 10333 37111
rect 10333 37077 10367 37111
rect 10367 37077 10376 37111
rect 10324 37068 10376 37077
rect 11888 37068 11940 37120
rect 12256 37111 12308 37120
rect 12256 37077 12265 37111
rect 12265 37077 12299 37111
rect 12299 37077 12308 37111
rect 12256 37068 12308 37077
rect 13544 37068 13596 37120
rect 15568 37068 15620 37120
rect 16672 37136 16724 37188
rect 17960 37247 18012 37256
rect 17960 37213 17969 37247
rect 17969 37213 18003 37247
rect 18003 37213 18012 37247
rect 18144 37247 18196 37256
rect 17960 37204 18012 37213
rect 18144 37213 18153 37247
rect 18153 37213 18187 37247
rect 18187 37213 18196 37247
rect 18144 37204 18196 37213
rect 18236 37247 18288 37256
rect 18236 37213 18245 37247
rect 18245 37213 18279 37247
rect 18279 37213 18288 37247
rect 18236 37204 18288 37213
rect 18604 37204 18656 37256
rect 20996 37204 21048 37256
rect 22192 37204 22244 37256
rect 25044 37204 25096 37256
rect 28908 37281 28917 37315
rect 28917 37281 28951 37315
rect 28951 37281 28960 37315
rect 28908 37272 28960 37281
rect 27252 37247 27304 37256
rect 27252 37213 27261 37247
rect 27261 37213 27295 37247
rect 27295 37213 27304 37247
rect 27252 37204 27304 37213
rect 18328 37136 18380 37188
rect 18420 37136 18472 37188
rect 21088 37179 21140 37188
rect 21088 37145 21097 37179
rect 21097 37145 21131 37179
rect 21131 37145 21140 37179
rect 21088 37136 21140 37145
rect 22100 37136 22152 37188
rect 25320 37136 25372 37188
rect 27620 37136 27672 37188
rect 19156 37068 19208 37120
rect 19340 37068 19392 37120
rect 20168 37068 20220 37120
rect 20720 37068 20772 37120
rect 23756 37068 23808 37120
rect 24492 37068 24544 37120
rect 26792 37111 26844 37120
rect 26792 37077 26801 37111
rect 26801 37077 26835 37111
rect 26835 37077 26844 37111
rect 26792 37068 26844 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 11888 36907 11940 36916
rect 11888 36873 11897 36907
rect 11897 36873 11931 36907
rect 11931 36873 11940 36907
rect 11888 36864 11940 36873
rect 13728 36864 13780 36916
rect 14096 36907 14148 36916
rect 14096 36873 14105 36907
rect 14105 36873 14139 36907
rect 14139 36873 14148 36907
rect 14096 36864 14148 36873
rect 16672 36864 16724 36916
rect 18696 36907 18748 36916
rect 18696 36873 18705 36907
rect 18705 36873 18739 36907
rect 18739 36873 18748 36907
rect 18696 36864 18748 36873
rect 8944 36728 8996 36780
rect 9864 36771 9916 36780
rect 9864 36737 9898 36771
rect 9898 36737 9916 36771
rect 9864 36728 9916 36737
rect 12532 36771 12584 36780
rect 12532 36737 12541 36771
rect 12541 36737 12575 36771
rect 12575 36737 12584 36771
rect 12532 36728 12584 36737
rect 16212 36796 16264 36848
rect 15568 36771 15620 36780
rect 12808 36660 12860 36712
rect 13820 36660 13872 36712
rect 11980 36592 12032 36644
rect 15568 36737 15577 36771
rect 15577 36737 15611 36771
rect 15611 36737 15620 36771
rect 15568 36728 15620 36737
rect 16948 36796 17000 36848
rect 19156 36839 19208 36848
rect 19156 36805 19165 36839
rect 19165 36805 19199 36839
rect 19199 36805 19208 36839
rect 19156 36796 19208 36805
rect 17684 36728 17736 36780
rect 16028 36660 16080 36712
rect 17592 36660 17644 36712
rect 17960 36660 18012 36712
rect 18328 36660 18380 36712
rect 19892 36728 19944 36780
rect 22376 36864 22428 36916
rect 23296 36864 23348 36916
rect 23756 36907 23808 36916
rect 23756 36873 23765 36907
rect 23765 36873 23799 36907
rect 23799 36873 23808 36907
rect 23756 36864 23808 36873
rect 26424 36907 26476 36916
rect 26424 36873 26433 36907
rect 26433 36873 26467 36907
rect 26467 36873 26476 36907
rect 26424 36864 26476 36873
rect 27620 36907 27672 36916
rect 27620 36873 27629 36907
rect 27629 36873 27663 36907
rect 27663 36873 27672 36907
rect 27620 36864 27672 36873
rect 20720 36771 20772 36780
rect 20720 36737 20729 36771
rect 20729 36737 20763 36771
rect 20763 36737 20772 36771
rect 26792 36796 26844 36848
rect 20720 36728 20772 36737
rect 20996 36660 21048 36712
rect 21088 36660 21140 36712
rect 22192 36771 22244 36780
rect 22192 36737 22201 36771
rect 22201 36737 22235 36771
rect 22235 36737 22244 36771
rect 22192 36728 22244 36737
rect 23388 36728 23440 36780
rect 23664 36771 23716 36780
rect 23664 36737 23673 36771
rect 23673 36737 23707 36771
rect 23707 36737 23716 36771
rect 23664 36728 23716 36737
rect 24492 36771 24544 36780
rect 24492 36737 24501 36771
rect 24501 36737 24535 36771
rect 24535 36737 24544 36771
rect 24492 36728 24544 36737
rect 25044 36771 25096 36780
rect 25044 36737 25053 36771
rect 25053 36737 25087 36771
rect 25087 36737 25096 36771
rect 25044 36728 25096 36737
rect 26332 36728 26384 36780
rect 19248 36592 19300 36644
rect 11152 36524 11204 36576
rect 11704 36524 11756 36576
rect 15844 36524 15896 36576
rect 19616 36524 19668 36576
rect 20168 36567 20220 36576
rect 20168 36533 20177 36567
rect 20177 36533 20211 36567
rect 20211 36533 20220 36567
rect 20168 36524 20220 36533
rect 21364 36524 21416 36576
rect 23664 36592 23716 36644
rect 24308 36567 24360 36576
rect 24308 36533 24317 36567
rect 24317 36533 24351 36567
rect 24351 36533 24360 36567
rect 24308 36524 24360 36533
rect 29828 36864 29880 36916
rect 28632 36839 28684 36848
rect 28632 36805 28641 36839
rect 28641 36805 28675 36839
rect 28675 36805 28684 36839
rect 28632 36796 28684 36805
rect 28540 36660 28592 36712
rect 29552 36524 29604 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 13176 36363 13228 36372
rect 13176 36329 13185 36363
rect 13185 36329 13219 36363
rect 13219 36329 13228 36363
rect 13176 36320 13228 36329
rect 16212 36363 16264 36372
rect 16212 36329 16221 36363
rect 16221 36329 16255 36363
rect 16255 36329 16264 36363
rect 16212 36320 16264 36329
rect 16948 36363 17000 36372
rect 16948 36329 16957 36363
rect 16957 36329 16991 36363
rect 16991 36329 17000 36363
rect 16948 36320 17000 36329
rect 18144 36320 18196 36372
rect 19616 36363 19668 36372
rect 19616 36329 19625 36363
rect 19625 36329 19659 36363
rect 19659 36329 19668 36363
rect 19616 36320 19668 36329
rect 19892 36252 19944 36304
rect 18420 36184 18472 36236
rect 19156 36184 19208 36236
rect 13084 36116 13136 36168
rect 16028 36116 16080 36168
rect 17684 36116 17736 36168
rect 19248 36159 19300 36168
rect 19248 36125 19257 36159
rect 19257 36125 19291 36159
rect 19291 36125 19300 36159
rect 19248 36116 19300 36125
rect 15568 36048 15620 36100
rect 17776 36048 17828 36100
rect 20628 36048 20680 36100
rect 22560 36252 22612 36304
rect 22100 36184 22152 36236
rect 37280 36320 37332 36372
rect 26332 36295 26384 36304
rect 26332 36261 26341 36295
rect 26341 36261 26375 36295
rect 26375 36261 26384 36295
rect 26332 36252 26384 36261
rect 29920 36252 29972 36304
rect 28540 36227 28592 36236
rect 28540 36193 28549 36227
rect 28549 36193 28583 36227
rect 28583 36193 28592 36227
rect 28540 36184 28592 36193
rect 21364 36159 21416 36168
rect 21364 36125 21373 36159
rect 21373 36125 21407 36159
rect 21407 36125 21416 36159
rect 26516 36159 26568 36168
rect 21364 36116 21416 36125
rect 26516 36125 26525 36159
rect 26525 36125 26559 36159
rect 26559 36125 26568 36159
rect 26516 36116 26568 36125
rect 28448 36159 28500 36168
rect 28448 36125 28457 36159
rect 28457 36125 28491 36159
rect 28491 36125 28500 36159
rect 28448 36116 28500 36125
rect 28816 36116 28868 36168
rect 22560 36048 22612 36100
rect 22928 36048 22980 36100
rect 25504 36091 25556 36100
rect 25504 36057 25513 36091
rect 25513 36057 25547 36091
rect 25547 36057 25556 36091
rect 25504 36048 25556 36057
rect 27896 36048 27948 36100
rect 11612 36023 11664 36032
rect 11612 35989 11621 36023
rect 11621 35989 11655 36023
rect 11655 35989 11664 36023
rect 11612 35980 11664 35989
rect 21364 35980 21416 36032
rect 22192 35980 22244 36032
rect 22468 36023 22520 36032
rect 22468 35989 22477 36023
rect 22477 35989 22511 36023
rect 22511 35989 22520 36023
rect 22468 35980 22520 35989
rect 25688 36023 25740 36032
rect 25688 35989 25713 36023
rect 25713 35989 25740 36023
rect 25872 36023 25924 36032
rect 25688 35980 25740 35989
rect 25872 35989 25881 36023
rect 25881 35989 25915 36023
rect 25915 35989 25924 36023
rect 25872 35980 25924 35989
rect 25964 35980 26016 36032
rect 28540 35980 28592 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 12992 35776 13044 35828
rect 14280 35776 14332 35828
rect 15108 35776 15160 35828
rect 15752 35776 15804 35828
rect 16672 35776 16724 35828
rect 17132 35776 17184 35828
rect 10324 35708 10376 35760
rect 10968 35640 11020 35692
rect 12440 35708 12492 35760
rect 12900 35708 12952 35760
rect 11612 35640 11664 35692
rect 15476 35683 15528 35692
rect 15476 35649 15485 35683
rect 15485 35649 15519 35683
rect 15519 35649 15528 35683
rect 15476 35640 15528 35649
rect 15752 35683 15804 35692
rect 12992 35572 13044 35624
rect 15752 35649 15761 35683
rect 15761 35649 15795 35683
rect 15795 35649 15804 35683
rect 15752 35640 15804 35649
rect 15844 35683 15896 35692
rect 15844 35649 15853 35683
rect 15853 35649 15887 35683
rect 15887 35649 15896 35683
rect 16672 35683 16724 35692
rect 15844 35640 15896 35649
rect 16672 35649 16681 35683
rect 16681 35649 16715 35683
rect 16715 35649 16724 35683
rect 16672 35640 16724 35649
rect 21916 35708 21968 35760
rect 22744 35708 22796 35760
rect 19156 35640 19208 35692
rect 19708 35615 19760 35624
rect 19708 35581 19717 35615
rect 19717 35581 19751 35615
rect 19751 35581 19760 35615
rect 19708 35572 19760 35581
rect 20076 35640 20128 35692
rect 21456 35640 21508 35692
rect 20628 35615 20680 35624
rect 20628 35581 20637 35615
rect 20637 35581 20671 35615
rect 20671 35581 20680 35615
rect 20628 35572 20680 35581
rect 15476 35504 15528 35556
rect 15660 35504 15712 35556
rect 22928 35640 22980 35692
rect 25044 35708 25096 35760
rect 25780 35708 25832 35760
rect 24308 35640 24360 35692
rect 26516 35776 26568 35828
rect 28264 35776 28316 35828
rect 28632 35776 28684 35828
rect 27896 35751 27948 35760
rect 27896 35717 27905 35751
rect 27905 35717 27939 35751
rect 27939 35717 27948 35751
rect 27896 35708 27948 35717
rect 28448 35640 28500 35692
rect 28724 35683 28776 35692
rect 28724 35649 28733 35683
rect 28733 35649 28767 35683
rect 28767 35649 28776 35683
rect 28724 35640 28776 35649
rect 28816 35640 28868 35692
rect 29736 35640 29788 35692
rect 22468 35572 22520 35624
rect 21640 35504 21692 35556
rect 25504 35547 25556 35556
rect 9956 35436 10008 35488
rect 12256 35436 12308 35488
rect 14004 35436 14056 35488
rect 16948 35436 17000 35488
rect 20996 35436 21048 35488
rect 25504 35513 25513 35547
rect 25513 35513 25547 35547
rect 25547 35513 25556 35547
rect 25504 35504 25556 35513
rect 22468 35479 22520 35488
rect 22468 35445 22477 35479
rect 22477 35445 22511 35479
rect 22511 35445 22520 35479
rect 22468 35436 22520 35445
rect 24492 35479 24544 35488
rect 24492 35445 24501 35479
rect 24501 35445 24535 35479
rect 24535 35445 24544 35479
rect 24492 35436 24544 35445
rect 25872 35479 25924 35488
rect 25872 35445 25881 35479
rect 25881 35445 25915 35479
rect 25915 35445 25924 35479
rect 25872 35436 25924 35445
rect 28172 35504 28224 35556
rect 28540 35504 28592 35556
rect 30564 35751 30616 35760
rect 30564 35717 30589 35751
rect 30589 35717 30616 35751
rect 30564 35708 30616 35717
rect 30840 35640 30892 35692
rect 37556 35572 37608 35624
rect 32128 35504 32180 35556
rect 30748 35479 30800 35488
rect 30748 35445 30757 35479
rect 30757 35445 30791 35479
rect 30791 35445 30800 35479
rect 30748 35436 30800 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 9864 35275 9916 35284
rect 9864 35241 9873 35275
rect 9873 35241 9907 35275
rect 9907 35241 9916 35275
rect 9864 35232 9916 35241
rect 11796 35275 11848 35284
rect 11796 35241 11805 35275
rect 11805 35241 11839 35275
rect 11839 35241 11848 35275
rect 11796 35232 11848 35241
rect 9864 35096 9916 35148
rect 10508 35071 10560 35080
rect 10508 35037 10517 35071
rect 10517 35037 10551 35071
rect 10551 35037 10560 35071
rect 10508 35028 10560 35037
rect 10968 35071 11020 35080
rect 10968 35037 10977 35071
rect 10977 35037 11011 35071
rect 11011 35037 11020 35071
rect 10968 35028 11020 35037
rect 11152 35071 11204 35080
rect 11152 35037 11161 35071
rect 11161 35037 11195 35071
rect 11195 35037 11204 35071
rect 11152 35028 11204 35037
rect 14096 35232 14148 35284
rect 12716 35207 12768 35216
rect 12716 35173 12725 35207
rect 12725 35173 12759 35207
rect 12759 35173 12768 35207
rect 12716 35164 12768 35173
rect 14464 35164 14516 35216
rect 15752 35232 15804 35284
rect 17960 35275 18012 35284
rect 17960 35241 17969 35275
rect 17969 35241 18003 35275
rect 18003 35241 18012 35275
rect 17960 35232 18012 35241
rect 19248 35275 19300 35284
rect 19248 35241 19257 35275
rect 19257 35241 19291 35275
rect 19291 35241 19300 35275
rect 19248 35232 19300 35241
rect 21732 35232 21784 35284
rect 21916 35232 21968 35284
rect 28172 35275 28224 35284
rect 12900 35028 12952 35080
rect 13176 35028 13228 35080
rect 14188 35071 14240 35080
rect 14188 35037 14198 35071
rect 14198 35037 14232 35071
rect 14232 35037 14240 35071
rect 14188 35028 14240 35037
rect 14648 35028 14700 35080
rect 15384 35028 15436 35080
rect 16488 35164 16540 35216
rect 21640 35207 21692 35216
rect 16212 35096 16264 35148
rect 19156 35096 19208 35148
rect 17684 35028 17736 35080
rect 12440 34960 12492 35012
rect 12992 34960 13044 35012
rect 14372 35003 14424 35012
rect 14372 34969 14381 35003
rect 14381 34969 14415 35003
rect 14415 34969 14424 35003
rect 14372 34960 14424 34969
rect 14924 34960 14976 35012
rect 18420 35028 18472 35080
rect 18880 34960 18932 35012
rect 19156 34960 19208 35012
rect 14556 34892 14608 34944
rect 15660 34892 15712 34944
rect 21640 35173 21649 35207
rect 21649 35173 21683 35207
rect 21683 35173 21692 35207
rect 21640 35164 21692 35173
rect 19708 35096 19760 35148
rect 20352 35028 20404 35080
rect 20628 35028 20680 35080
rect 20996 35028 21048 35080
rect 22192 35096 22244 35148
rect 28172 35241 28181 35275
rect 28181 35241 28215 35275
rect 28215 35241 28224 35275
rect 28172 35232 28224 35241
rect 30380 35275 30432 35284
rect 30380 35241 30389 35275
rect 30389 35241 30423 35275
rect 30423 35241 30432 35275
rect 30380 35232 30432 35241
rect 31024 35275 31076 35284
rect 31024 35241 31033 35275
rect 31033 35241 31067 35275
rect 31067 35241 31076 35275
rect 31024 35232 31076 35241
rect 25504 35164 25556 35216
rect 30196 35207 30248 35216
rect 30196 35173 30205 35207
rect 30205 35173 30239 35207
rect 30239 35173 30248 35207
rect 30196 35164 30248 35173
rect 30472 35164 30524 35216
rect 32404 35096 32456 35148
rect 22468 35071 22520 35080
rect 22468 35037 22477 35071
rect 22477 35037 22511 35071
rect 22511 35037 22520 35071
rect 22468 35028 22520 35037
rect 25964 35071 26016 35080
rect 25964 35037 25973 35071
rect 25973 35037 26007 35071
rect 26007 35037 26016 35071
rect 25964 35028 26016 35037
rect 26332 35028 26384 35080
rect 27804 35071 27856 35080
rect 27804 35037 27813 35071
rect 27813 35037 27847 35071
rect 27847 35037 27856 35071
rect 27804 35028 27856 35037
rect 28540 35028 28592 35080
rect 29092 35028 29144 35080
rect 30564 35028 30616 35080
rect 31116 35028 31168 35080
rect 22560 34960 22612 35012
rect 23940 34960 23992 35012
rect 25688 34960 25740 35012
rect 30840 35003 30892 35012
rect 30840 34969 30849 35003
rect 30849 34969 30883 35003
rect 30883 34969 30892 35003
rect 30840 34960 30892 34969
rect 23572 34892 23624 34944
rect 23848 34935 23900 34944
rect 23848 34901 23857 34935
rect 23857 34901 23891 34935
rect 23891 34901 23900 34935
rect 23848 34892 23900 34901
rect 25320 34892 25372 34944
rect 28080 34892 28132 34944
rect 30380 34892 30432 34944
rect 31576 34892 31628 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 9588 34688 9640 34740
rect 12624 34688 12676 34740
rect 13728 34688 13780 34740
rect 13912 34688 13964 34740
rect 8944 34595 8996 34604
rect 8944 34561 8953 34595
rect 8953 34561 8987 34595
rect 8987 34561 8996 34595
rect 8944 34552 8996 34561
rect 10416 34620 10468 34672
rect 12900 34620 12952 34672
rect 12072 34595 12124 34604
rect 9772 34527 9824 34536
rect 9772 34493 9781 34527
rect 9781 34493 9815 34527
rect 9815 34493 9824 34527
rect 9772 34484 9824 34493
rect 12072 34561 12081 34595
rect 12081 34561 12115 34595
rect 12115 34561 12124 34595
rect 12072 34552 12124 34561
rect 12256 34595 12308 34604
rect 12256 34561 12263 34595
rect 12263 34561 12308 34595
rect 12256 34552 12308 34561
rect 10232 34484 10284 34536
rect 10508 34484 10560 34536
rect 12624 34552 12676 34604
rect 13636 34595 13688 34604
rect 13636 34561 13645 34595
rect 13645 34561 13679 34595
rect 13679 34561 13688 34595
rect 13636 34552 13688 34561
rect 16488 34620 16540 34672
rect 14648 34552 14700 34604
rect 15108 34552 15160 34604
rect 9864 34416 9916 34468
rect 14280 34484 14332 34536
rect 17776 34688 17828 34740
rect 17868 34620 17920 34672
rect 17960 34620 18012 34672
rect 18972 34663 19024 34672
rect 18972 34629 18981 34663
rect 18981 34629 19015 34663
rect 19015 34629 19024 34663
rect 18972 34620 19024 34629
rect 19340 34688 19392 34740
rect 19156 34663 19208 34672
rect 19156 34629 19191 34663
rect 19191 34629 19208 34663
rect 19156 34620 19208 34629
rect 19708 34620 19760 34672
rect 16856 34595 16908 34604
rect 16856 34561 16865 34595
rect 16865 34561 16899 34595
rect 16899 34561 16908 34595
rect 16856 34552 16908 34561
rect 14372 34416 14424 34468
rect 17132 34595 17184 34604
rect 17132 34561 17167 34595
rect 17167 34561 17184 34595
rect 17132 34552 17184 34561
rect 18328 34552 18380 34604
rect 20904 34688 20956 34740
rect 21640 34688 21692 34740
rect 22100 34688 22152 34740
rect 22744 34731 22796 34740
rect 22744 34697 22753 34731
rect 22753 34697 22787 34731
rect 22787 34697 22796 34731
rect 22744 34688 22796 34697
rect 24216 34688 24268 34740
rect 25780 34731 25832 34740
rect 25780 34697 25789 34731
rect 25789 34697 25823 34731
rect 25823 34697 25832 34731
rect 25780 34688 25832 34697
rect 27988 34731 28040 34740
rect 27988 34697 27997 34731
rect 27997 34697 28031 34731
rect 28031 34697 28040 34731
rect 27988 34688 28040 34697
rect 29736 34731 29788 34740
rect 29736 34697 29745 34731
rect 29745 34697 29779 34731
rect 29779 34697 29788 34731
rect 29736 34688 29788 34697
rect 20352 34620 20404 34672
rect 21456 34620 21508 34672
rect 21824 34620 21876 34672
rect 17960 34416 18012 34468
rect 16672 34391 16724 34400
rect 16672 34357 16681 34391
rect 16681 34357 16715 34391
rect 16715 34357 16724 34391
rect 16672 34348 16724 34357
rect 16856 34348 16908 34400
rect 19340 34527 19392 34536
rect 19340 34493 19349 34527
rect 19349 34493 19383 34527
rect 19383 34493 19392 34527
rect 19340 34484 19392 34493
rect 20352 34484 20404 34536
rect 21824 34527 21876 34536
rect 18972 34416 19024 34468
rect 19708 34416 19760 34468
rect 21824 34493 21833 34527
rect 21833 34493 21867 34527
rect 21867 34493 21876 34527
rect 21824 34484 21876 34493
rect 22100 34552 22152 34604
rect 23572 34620 23624 34672
rect 20904 34416 20956 34468
rect 22100 34416 22152 34468
rect 23940 34484 23992 34536
rect 26332 34552 26384 34604
rect 28540 34552 28592 34604
rect 25964 34484 26016 34536
rect 26148 34484 26200 34536
rect 28264 34484 28316 34536
rect 28908 34552 28960 34604
rect 30288 34552 30340 34604
rect 31208 34552 31260 34604
rect 29092 34484 29144 34536
rect 22836 34416 22888 34468
rect 23296 34416 23348 34468
rect 27804 34459 27856 34468
rect 27804 34425 27813 34459
rect 27813 34425 27847 34459
rect 27847 34425 27856 34459
rect 27804 34416 27856 34425
rect 29644 34459 29696 34468
rect 29644 34425 29653 34459
rect 29653 34425 29687 34459
rect 29687 34425 29696 34459
rect 29644 34416 29696 34425
rect 18604 34348 18656 34400
rect 19248 34348 19300 34400
rect 20444 34348 20496 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 9404 34187 9456 34196
rect 9404 34153 9413 34187
rect 9413 34153 9447 34187
rect 9447 34153 9456 34187
rect 9404 34144 9456 34153
rect 10692 34144 10744 34196
rect 14464 34144 14516 34196
rect 15476 34144 15528 34196
rect 19432 34144 19484 34196
rect 20536 34144 20588 34196
rect 23848 34144 23900 34196
rect 30748 34144 30800 34196
rect 31208 34187 31260 34196
rect 31208 34153 31217 34187
rect 31217 34153 31251 34187
rect 31251 34153 31260 34187
rect 31208 34144 31260 34153
rect 9864 34076 9916 34128
rect 10968 34076 11020 34128
rect 9956 33940 10008 33992
rect 10232 33940 10284 33992
rect 10692 33940 10744 33992
rect 11980 33940 12032 33992
rect 12348 33983 12400 33992
rect 12348 33949 12355 33983
rect 12355 33949 12400 33983
rect 12348 33940 12400 33949
rect 14464 34008 14516 34060
rect 12624 33940 12676 33992
rect 11520 33872 11572 33924
rect 13084 33872 13136 33924
rect 13360 33940 13412 33992
rect 16672 34076 16724 34128
rect 18236 34076 18288 34128
rect 16488 33983 16540 33992
rect 12624 33804 12676 33856
rect 13820 33804 13872 33856
rect 14280 33804 14332 33856
rect 15568 33872 15620 33924
rect 16488 33949 16497 33983
rect 16497 33949 16531 33983
rect 16531 33949 16540 33983
rect 16488 33940 16540 33949
rect 16764 34008 16816 34060
rect 16672 33983 16724 33992
rect 16672 33949 16686 33983
rect 16686 33949 16720 33983
rect 16720 33949 16724 33983
rect 17408 33983 17460 33992
rect 16672 33940 16724 33949
rect 17408 33949 17417 33983
rect 17417 33949 17451 33983
rect 17451 33949 17460 33983
rect 17408 33940 17460 33949
rect 17960 33940 18012 33992
rect 19248 33983 19300 33992
rect 19248 33949 19257 33983
rect 19257 33949 19291 33983
rect 19291 33949 19300 33983
rect 19248 33940 19300 33949
rect 19432 33983 19484 33992
rect 19432 33949 19439 33983
rect 19439 33949 19484 33983
rect 19432 33940 19484 33949
rect 20076 34008 20128 34060
rect 20720 34008 20772 34060
rect 30196 34119 30248 34128
rect 30196 34085 30205 34119
rect 30205 34085 30239 34119
rect 30239 34085 30248 34119
rect 30196 34076 30248 34085
rect 16948 33872 17000 33924
rect 17868 33872 17920 33924
rect 19064 33872 19116 33924
rect 19624 33915 19676 33924
rect 19624 33881 19645 33915
rect 19645 33881 19676 33915
rect 20444 33983 20496 33992
rect 20444 33949 20453 33983
rect 20453 33949 20487 33983
rect 20487 33949 20496 33983
rect 20444 33940 20496 33949
rect 20536 33983 20588 33992
rect 20536 33949 20546 33983
rect 20546 33949 20580 33983
rect 20580 33949 20588 33983
rect 20536 33940 20588 33949
rect 21640 33983 21692 33992
rect 21640 33949 21649 33983
rect 21649 33949 21683 33983
rect 21683 33949 21692 33983
rect 21640 33940 21692 33949
rect 21824 33983 21876 33992
rect 21824 33949 21831 33983
rect 21831 33949 21876 33983
rect 21824 33940 21876 33949
rect 22008 33983 22060 33992
rect 22008 33949 22017 33983
rect 22017 33949 22051 33983
rect 22051 33949 22060 33983
rect 22008 33940 22060 33949
rect 23296 33983 23348 33992
rect 23296 33949 23305 33983
rect 23305 33949 23339 33983
rect 23339 33949 23348 33983
rect 23296 33940 23348 33949
rect 19624 33872 19676 33881
rect 15108 33804 15160 33856
rect 16672 33804 16724 33856
rect 17316 33804 17368 33856
rect 18236 33804 18288 33856
rect 19984 33804 20036 33856
rect 21088 33847 21140 33856
rect 21088 33813 21097 33847
rect 21097 33813 21131 33847
rect 21131 33813 21140 33847
rect 21088 33804 21140 33813
rect 22468 33804 22520 33856
rect 23664 33847 23716 33856
rect 23664 33813 23673 33847
rect 23673 33813 23707 33847
rect 23707 33813 23716 33847
rect 23664 33804 23716 33813
rect 28080 33983 28132 33992
rect 28080 33949 28089 33983
rect 28089 33949 28123 33983
rect 28123 33949 28132 33983
rect 28080 33940 28132 33949
rect 29552 33983 29604 33992
rect 29552 33949 29561 33983
rect 29561 33949 29595 33983
rect 29595 33949 29604 33983
rect 29552 33940 29604 33949
rect 30564 33940 30616 33992
rect 24768 33872 24820 33924
rect 26516 33872 26568 33924
rect 24032 33804 24084 33856
rect 25044 33804 25096 33856
rect 27528 33804 27580 33856
rect 27896 33847 27948 33856
rect 27896 33813 27905 33847
rect 27905 33813 27939 33847
rect 27939 33813 27948 33847
rect 27896 33804 27948 33813
rect 30288 33804 30340 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 10416 33643 10468 33652
rect 10416 33609 10425 33643
rect 10425 33609 10459 33643
rect 10459 33609 10468 33643
rect 10416 33600 10468 33609
rect 11980 33643 12032 33652
rect 11980 33609 11989 33643
rect 11989 33609 12023 33643
rect 12023 33609 12032 33643
rect 11980 33600 12032 33609
rect 12164 33600 12216 33652
rect 13636 33643 13688 33652
rect 10784 33532 10836 33584
rect 10968 33532 11020 33584
rect 11060 33532 11112 33584
rect 13636 33609 13645 33643
rect 13645 33609 13679 33643
rect 13679 33609 13688 33643
rect 13636 33600 13688 33609
rect 12440 33575 12492 33584
rect 12440 33541 12475 33575
rect 12475 33541 12492 33575
rect 12440 33532 12492 33541
rect 13544 33532 13596 33584
rect 16488 33600 16540 33652
rect 17868 33600 17920 33652
rect 18328 33600 18380 33652
rect 18696 33600 18748 33652
rect 20444 33600 20496 33652
rect 21640 33600 21692 33652
rect 23296 33600 23348 33652
rect 14280 33532 14332 33584
rect 10600 33464 10652 33516
rect 12164 33507 12216 33516
rect 12164 33473 12173 33507
rect 12173 33473 12207 33507
rect 12207 33473 12216 33507
rect 12164 33464 12216 33473
rect 13636 33464 13688 33516
rect 14832 33532 14884 33584
rect 15384 33532 15436 33584
rect 16948 33532 17000 33584
rect 17132 33532 17184 33584
rect 18972 33532 19024 33584
rect 21548 33532 21600 33584
rect 21824 33532 21876 33584
rect 26516 33600 26568 33652
rect 27252 33600 27304 33652
rect 30380 33600 30432 33652
rect 27896 33532 27948 33584
rect 30288 33575 30340 33584
rect 30288 33541 30297 33575
rect 30297 33541 30331 33575
rect 30331 33541 30340 33575
rect 30288 33532 30340 33541
rect 14924 33507 14976 33516
rect 12348 33396 12400 33448
rect 12716 33396 12768 33448
rect 14924 33473 14933 33507
rect 14933 33473 14967 33507
rect 14967 33473 14976 33507
rect 14924 33464 14976 33473
rect 15844 33507 15896 33516
rect 14832 33396 14884 33448
rect 14924 33328 14976 33380
rect 15016 33328 15068 33380
rect 15844 33473 15853 33507
rect 15853 33473 15887 33507
rect 15887 33473 15896 33507
rect 15844 33464 15896 33473
rect 18144 33464 18196 33516
rect 18236 33507 18288 33516
rect 18236 33473 18245 33507
rect 18245 33473 18279 33507
rect 18279 33473 18288 33507
rect 18236 33464 18288 33473
rect 18604 33464 18656 33516
rect 20996 33507 21048 33516
rect 20996 33473 21031 33507
rect 21031 33473 21048 33507
rect 20996 33464 21048 33473
rect 22284 33464 22336 33516
rect 24124 33507 24176 33516
rect 24124 33473 24133 33507
rect 24133 33473 24167 33507
rect 24167 33473 24176 33507
rect 24124 33464 24176 33473
rect 24584 33464 24636 33516
rect 25044 33507 25096 33516
rect 25044 33473 25053 33507
rect 25053 33473 25087 33507
rect 25087 33473 25096 33507
rect 25044 33464 25096 33473
rect 27528 33507 27580 33516
rect 27528 33473 27537 33507
rect 27537 33473 27571 33507
rect 27571 33473 27580 33507
rect 27528 33464 27580 33473
rect 27804 33507 27856 33516
rect 27804 33473 27838 33507
rect 27838 33473 27856 33507
rect 27804 33464 27856 33473
rect 29000 33464 29052 33516
rect 29552 33464 29604 33516
rect 30564 33464 30616 33516
rect 30840 33464 30892 33516
rect 14280 33260 14332 33312
rect 14648 33260 14700 33312
rect 14832 33260 14884 33312
rect 16212 33396 16264 33448
rect 16672 33439 16724 33448
rect 16672 33405 16681 33439
rect 16681 33405 16715 33439
rect 16715 33405 16724 33439
rect 16672 33396 16724 33405
rect 16856 33396 16908 33448
rect 17776 33396 17828 33448
rect 18052 33396 18104 33448
rect 20352 33396 20404 33448
rect 20444 33396 20496 33448
rect 20904 33396 20956 33448
rect 22192 33439 22244 33448
rect 22192 33405 22201 33439
rect 22201 33405 22235 33439
rect 22235 33405 22244 33439
rect 22192 33396 22244 33405
rect 23480 33260 23532 33312
rect 28540 33260 28592 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 18328 33056 18380 33108
rect 19340 33056 19392 33108
rect 20076 33056 20128 33108
rect 22284 33056 22336 33108
rect 28724 33056 28776 33108
rect 9956 32988 10008 33040
rect 12072 33031 12124 33040
rect 12072 32997 12081 33031
rect 12081 32997 12115 33031
rect 12115 32997 12124 33031
rect 12072 32988 12124 32997
rect 13268 32988 13320 33040
rect 12164 32920 12216 32972
rect 9496 32784 9548 32836
rect 9680 32759 9732 32768
rect 9680 32725 9689 32759
rect 9689 32725 9723 32759
rect 9723 32725 9732 32759
rect 9680 32716 9732 32725
rect 10232 32852 10284 32904
rect 10784 32895 10836 32904
rect 10784 32861 10793 32895
rect 10793 32861 10827 32895
rect 10827 32861 10836 32895
rect 10784 32852 10836 32861
rect 11060 32852 11112 32904
rect 13636 32920 13688 32972
rect 15568 32988 15620 33040
rect 12348 32895 12400 32904
rect 12348 32861 12357 32895
rect 12357 32861 12391 32895
rect 12391 32861 12400 32895
rect 12716 32895 12768 32904
rect 12348 32852 12400 32861
rect 12716 32861 12725 32895
rect 12725 32861 12759 32895
rect 12759 32861 12768 32895
rect 12716 32852 12768 32861
rect 13360 32852 13412 32904
rect 17408 32920 17460 32972
rect 14188 32852 14240 32904
rect 14924 32852 14976 32904
rect 15660 32852 15712 32904
rect 20536 32988 20588 33040
rect 17868 32963 17920 32972
rect 17868 32929 17877 32963
rect 17877 32929 17911 32963
rect 17911 32929 17920 32963
rect 17868 32920 17920 32929
rect 18604 32852 18656 32904
rect 19248 32895 19300 32904
rect 19248 32861 19257 32895
rect 19257 32861 19291 32895
rect 19291 32861 19300 32895
rect 19248 32852 19300 32861
rect 19432 32895 19484 32904
rect 19432 32861 19441 32895
rect 19441 32861 19475 32895
rect 19475 32861 19484 32895
rect 19432 32852 19484 32861
rect 19524 32852 19576 32904
rect 19708 32895 19760 32904
rect 19708 32861 19717 32895
rect 19717 32861 19751 32895
rect 19751 32861 19760 32895
rect 19708 32852 19760 32861
rect 10600 32784 10652 32836
rect 11888 32716 11940 32768
rect 12808 32784 12860 32836
rect 18236 32784 18288 32836
rect 22100 32895 22152 32904
rect 22100 32861 22109 32895
rect 22109 32861 22143 32895
rect 22143 32861 22152 32895
rect 22100 32852 22152 32861
rect 22744 32852 22796 32904
rect 25044 32852 25096 32904
rect 27620 32895 27672 32904
rect 27620 32861 27629 32895
rect 27629 32861 27663 32895
rect 27663 32861 27672 32895
rect 27620 32852 27672 32861
rect 30656 32852 30708 32904
rect 14832 32716 14884 32768
rect 17684 32716 17736 32768
rect 20352 32716 20404 32768
rect 23296 32784 23348 32836
rect 23572 32827 23624 32836
rect 23572 32793 23581 32827
rect 23581 32793 23615 32827
rect 23615 32793 23624 32827
rect 23572 32784 23624 32793
rect 25320 32784 25372 32836
rect 28172 32784 28224 32836
rect 23480 32716 23532 32768
rect 26148 32716 26200 32768
rect 30564 32759 30616 32768
rect 30564 32725 30573 32759
rect 30573 32725 30607 32759
rect 30607 32725 30616 32759
rect 30564 32716 30616 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 11060 32512 11112 32564
rect 15384 32512 15436 32564
rect 20444 32555 20496 32564
rect 9680 32444 9732 32496
rect 10784 32444 10836 32496
rect 5908 32376 5960 32428
rect 8116 32376 8168 32428
rect 11704 32419 11756 32428
rect 11704 32385 11713 32419
rect 11713 32385 11747 32419
rect 11747 32385 11756 32419
rect 11704 32376 11756 32385
rect 13268 32376 13320 32428
rect 6736 32308 6788 32360
rect 9312 32308 9364 32360
rect 11980 32308 12032 32360
rect 13820 32308 13872 32360
rect 14464 32444 14516 32496
rect 15660 32444 15712 32496
rect 14648 32419 14700 32428
rect 14648 32385 14657 32419
rect 14657 32385 14691 32419
rect 14691 32385 14700 32419
rect 14648 32376 14700 32385
rect 14832 32419 14884 32428
rect 14832 32385 14839 32419
rect 14839 32385 14884 32419
rect 14832 32376 14884 32385
rect 15108 32419 15160 32428
rect 15108 32385 15122 32419
rect 15122 32385 15156 32419
rect 15156 32385 15160 32419
rect 15108 32376 15160 32385
rect 16764 32419 16816 32428
rect 15016 32308 15068 32360
rect 16764 32385 16773 32419
rect 16773 32385 16807 32419
rect 16807 32385 16816 32419
rect 16764 32376 16816 32385
rect 17868 32444 17920 32496
rect 19248 32444 19300 32496
rect 20444 32521 20453 32555
rect 20453 32521 20487 32555
rect 20487 32521 20496 32555
rect 20444 32512 20496 32521
rect 22100 32512 22152 32564
rect 22744 32512 22796 32564
rect 23296 32512 23348 32564
rect 23664 32512 23716 32564
rect 25320 32555 25372 32564
rect 25320 32521 25329 32555
rect 25329 32521 25363 32555
rect 25363 32521 25372 32555
rect 25320 32512 25372 32521
rect 25780 32512 25832 32564
rect 27712 32512 27764 32564
rect 28172 32555 28224 32564
rect 28172 32521 28181 32555
rect 28181 32521 28215 32555
rect 28215 32521 28224 32555
rect 28172 32512 28224 32521
rect 28724 32512 28776 32564
rect 30564 32444 30616 32496
rect 17132 32419 17184 32428
rect 17132 32385 17141 32419
rect 17141 32385 17175 32419
rect 17175 32385 17184 32419
rect 17132 32376 17184 32385
rect 17316 32376 17368 32428
rect 20352 32419 20404 32428
rect 20352 32385 20361 32419
rect 20361 32385 20395 32419
rect 20395 32385 20404 32419
rect 20352 32376 20404 32385
rect 24124 32376 24176 32428
rect 24400 32419 24452 32428
rect 24400 32385 24409 32419
rect 24409 32385 24443 32419
rect 24443 32385 24452 32419
rect 24400 32376 24452 32385
rect 24584 32419 24636 32428
rect 24584 32385 24593 32419
rect 24593 32385 24627 32419
rect 24627 32385 24636 32419
rect 24584 32376 24636 32385
rect 25596 32376 25648 32428
rect 16672 32308 16724 32360
rect 17868 32308 17920 32360
rect 5264 32172 5316 32224
rect 6368 32215 6420 32224
rect 6368 32181 6377 32215
rect 6377 32181 6411 32215
rect 6411 32181 6420 32215
rect 6368 32172 6420 32181
rect 7748 32215 7800 32224
rect 7748 32181 7757 32215
rect 7757 32181 7791 32215
rect 7791 32181 7800 32215
rect 7748 32172 7800 32181
rect 9496 32172 9548 32224
rect 15200 32240 15252 32292
rect 15568 32240 15620 32292
rect 11060 32172 11112 32224
rect 13636 32215 13688 32224
rect 13636 32181 13645 32215
rect 13645 32181 13679 32215
rect 13679 32181 13688 32215
rect 13636 32172 13688 32181
rect 15384 32172 15436 32224
rect 16672 32172 16724 32224
rect 17500 32172 17552 32224
rect 20536 32308 20588 32360
rect 22100 32308 22152 32360
rect 19524 32240 19576 32292
rect 20444 32240 20496 32292
rect 25320 32308 25372 32360
rect 25780 32419 25832 32428
rect 25780 32385 25789 32419
rect 25789 32385 25823 32419
rect 25823 32385 25832 32419
rect 27436 32419 27488 32428
rect 25780 32376 25832 32385
rect 27436 32385 27445 32419
rect 27445 32385 27479 32419
rect 27479 32385 27488 32419
rect 27436 32376 27488 32385
rect 26148 32308 26200 32360
rect 25872 32240 25924 32292
rect 27712 32419 27764 32428
rect 27712 32385 27721 32419
rect 27721 32385 27755 32419
rect 27755 32385 27764 32419
rect 28356 32419 28408 32428
rect 27712 32376 27764 32385
rect 28356 32385 28365 32419
rect 28365 32385 28399 32419
rect 28399 32385 28408 32419
rect 28356 32376 28408 32385
rect 30196 32351 30248 32360
rect 30196 32317 30205 32351
rect 30205 32317 30239 32351
rect 30239 32317 30248 32351
rect 30196 32308 30248 32317
rect 28540 32240 28592 32292
rect 18236 32172 18288 32224
rect 24032 32172 24084 32224
rect 27804 32172 27856 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 11704 31968 11756 32020
rect 11980 31968 12032 32020
rect 13820 31968 13872 32020
rect 14188 31968 14240 32020
rect 15200 31968 15252 32020
rect 17316 31968 17368 32020
rect 17500 31968 17552 32020
rect 13636 31832 13688 31884
rect 4988 31807 5040 31816
rect 4988 31773 4997 31807
rect 4997 31773 5031 31807
rect 5031 31773 5040 31807
rect 7012 31807 7064 31816
rect 4988 31764 5040 31773
rect 5264 31739 5316 31748
rect 5264 31705 5298 31739
rect 5298 31705 5316 31739
rect 5264 31696 5316 31705
rect 7012 31773 7021 31807
rect 7021 31773 7055 31807
rect 7055 31773 7064 31807
rect 7012 31764 7064 31773
rect 7748 31764 7800 31816
rect 9036 31764 9088 31816
rect 9312 31764 9364 31816
rect 14740 31832 14792 31884
rect 16764 31900 16816 31952
rect 14648 31764 14700 31816
rect 15568 31764 15620 31816
rect 18052 31807 18104 31816
rect 18052 31773 18061 31807
rect 18061 31773 18095 31807
rect 18095 31773 18104 31807
rect 18052 31764 18104 31773
rect 18236 31900 18288 31952
rect 18788 31832 18840 31884
rect 19432 31968 19484 32020
rect 23572 31968 23624 32020
rect 24032 31968 24084 32020
rect 25596 31968 25648 32020
rect 27436 31968 27488 32020
rect 30472 32011 30524 32020
rect 30472 31977 30481 32011
rect 30481 31977 30515 32011
rect 30515 31977 30524 32011
rect 30472 31968 30524 31977
rect 30656 32011 30708 32020
rect 30656 31977 30665 32011
rect 30665 31977 30699 32011
rect 30699 31977 30708 32011
rect 30656 31968 30708 31977
rect 22008 31943 22060 31952
rect 22008 31909 22017 31943
rect 22017 31909 22051 31943
rect 22051 31909 22060 31943
rect 22008 31900 22060 31909
rect 29644 31900 29696 31952
rect 20536 31832 20588 31884
rect 6828 31696 6880 31748
rect 9588 31696 9640 31748
rect 17776 31696 17828 31748
rect 17960 31696 18012 31748
rect 6368 31671 6420 31680
rect 6368 31637 6377 31671
rect 6377 31637 6411 31671
rect 6411 31637 6420 31671
rect 6368 31628 6420 31637
rect 8392 31671 8444 31680
rect 8392 31637 8401 31671
rect 8401 31637 8435 31671
rect 8435 31637 8444 31671
rect 8392 31628 8444 31637
rect 8944 31628 8996 31680
rect 13636 31628 13688 31680
rect 18144 31628 18196 31680
rect 18696 31764 18748 31816
rect 19340 31764 19392 31816
rect 19432 31696 19484 31748
rect 20444 31764 20496 31816
rect 22192 31832 22244 31884
rect 25872 31875 25924 31884
rect 25872 31841 25881 31875
rect 25881 31841 25915 31875
rect 25915 31841 25924 31875
rect 25872 31832 25924 31841
rect 27804 31875 27856 31884
rect 27804 31841 27813 31875
rect 27813 31841 27847 31875
rect 27847 31841 27856 31875
rect 27804 31832 27856 31841
rect 20904 31739 20956 31748
rect 20904 31705 20938 31739
rect 20938 31705 20956 31739
rect 20904 31696 20956 31705
rect 21180 31696 21232 31748
rect 21732 31696 21784 31748
rect 22100 31696 22152 31748
rect 23112 31696 23164 31748
rect 24124 31696 24176 31748
rect 27988 31764 28040 31816
rect 30748 31764 30800 31816
rect 31300 31807 31352 31816
rect 31300 31773 31309 31807
rect 31309 31773 31343 31807
rect 31343 31773 31352 31807
rect 31300 31764 31352 31773
rect 23664 31628 23716 31680
rect 24400 31628 24452 31680
rect 25412 31671 25464 31680
rect 25412 31637 25421 31671
rect 25421 31637 25455 31671
rect 25455 31637 25464 31671
rect 25412 31628 25464 31637
rect 27528 31628 27580 31680
rect 30472 31671 30524 31680
rect 30472 31637 30481 31671
rect 30481 31637 30515 31671
rect 30515 31637 30524 31671
rect 30472 31628 30524 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 5908 31424 5960 31476
rect 6552 31467 6604 31476
rect 6552 31433 6577 31467
rect 6577 31433 6604 31467
rect 6736 31467 6788 31476
rect 6552 31424 6604 31433
rect 6736 31433 6745 31467
rect 6745 31433 6779 31467
rect 6779 31433 6788 31467
rect 6736 31424 6788 31433
rect 9588 31467 9640 31476
rect 9588 31433 9597 31467
rect 9597 31433 9631 31467
rect 9631 31433 9640 31467
rect 9588 31424 9640 31433
rect 9956 31424 10008 31476
rect 12808 31424 12860 31476
rect 13636 31424 13688 31476
rect 13820 31424 13872 31476
rect 14648 31424 14700 31476
rect 18236 31424 18288 31476
rect 20904 31424 20956 31476
rect 21180 31467 21232 31476
rect 21180 31433 21189 31467
rect 21189 31433 21223 31467
rect 21223 31433 21232 31467
rect 21180 31424 21232 31433
rect 21824 31467 21876 31476
rect 21824 31433 21833 31467
rect 21833 31433 21867 31467
rect 21867 31433 21876 31467
rect 27528 31467 27580 31476
rect 21824 31424 21876 31433
rect 6736 31288 6788 31340
rect 7012 31288 7064 31340
rect 7288 31288 7340 31340
rect 9680 31288 9732 31340
rect 10232 31331 10284 31340
rect 10232 31297 10241 31331
rect 10241 31297 10275 31331
rect 10275 31297 10284 31331
rect 10232 31288 10284 31297
rect 16488 31356 16540 31408
rect 18512 31356 18564 31408
rect 18696 31356 18748 31408
rect 19432 31356 19484 31408
rect 27528 31433 27537 31467
rect 27537 31433 27571 31467
rect 27571 31433 27580 31467
rect 27528 31424 27580 31433
rect 28356 31424 28408 31476
rect 30472 31424 30524 31476
rect 13544 31331 13596 31340
rect 13544 31297 13553 31331
rect 13553 31297 13587 31331
rect 13587 31297 13596 31331
rect 13544 31288 13596 31297
rect 13820 31331 13872 31340
rect 13820 31297 13829 31331
rect 13829 31297 13863 31331
rect 13863 31297 13872 31331
rect 13820 31288 13872 31297
rect 14188 31288 14240 31340
rect 14372 31288 14424 31340
rect 16856 31331 16908 31340
rect 16856 31297 16865 31331
rect 16865 31297 16899 31331
rect 16899 31297 16908 31331
rect 16856 31288 16908 31297
rect 17132 31288 17184 31340
rect 18144 31331 18196 31340
rect 18144 31297 18153 31331
rect 18153 31297 18187 31331
rect 18187 31297 18196 31331
rect 18144 31288 18196 31297
rect 20812 31288 20864 31340
rect 24216 31356 24268 31408
rect 11060 31220 11112 31272
rect 18236 31220 18288 31272
rect 22100 31288 22152 31340
rect 22284 31331 22336 31340
rect 22284 31297 22293 31331
rect 22293 31297 22327 31331
rect 22327 31297 22336 31331
rect 22284 31288 22336 31297
rect 22008 31220 22060 31272
rect 23572 31263 23624 31272
rect 23572 31229 23581 31263
rect 23581 31229 23615 31263
rect 23615 31229 23624 31263
rect 23572 31220 23624 31229
rect 18328 31195 18380 31204
rect 18328 31161 18337 31195
rect 18337 31161 18371 31195
rect 18371 31161 18380 31195
rect 29000 31356 29052 31408
rect 25044 31288 25096 31340
rect 25228 31331 25280 31340
rect 25228 31297 25262 31331
rect 25262 31297 25280 31331
rect 27988 31331 28040 31340
rect 25228 31288 25280 31297
rect 27988 31297 27997 31331
rect 27997 31297 28031 31331
rect 28031 31297 28040 31331
rect 27988 31288 28040 31297
rect 30104 31356 30156 31408
rect 29184 31331 29236 31340
rect 29184 31297 29218 31331
rect 29218 31297 29236 31331
rect 30748 31331 30800 31340
rect 29184 31288 29236 31297
rect 18328 31152 18380 31161
rect 27988 31152 28040 31204
rect 5632 31127 5684 31136
rect 5632 31093 5641 31127
rect 5641 31093 5675 31127
rect 5675 31093 5684 31127
rect 5632 31084 5684 31093
rect 6368 31084 6420 31136
rect 8576 31127 8628 31136
rect 8576 31093 8585 31127
rect 8585 31093 8619 31127
rect 8619 31093 8628 31127
rect 8576 31084 8628 31093
rect 15660 31127 15712 31136
rect 15660 31093 15669 31127
rect 15669 31093 15703 31127
rect 15703 31093 15712 31127
rect 15660 31084 15712 31093
rect 17132 31084 17184 31136
rect 17224 31084 17276 31136
rect 20352 31084 20404 31136
rect 23296 31084 23348 31136
rect 26148 31084 26200 31136
rect 28632 31084 28684 31136
rect 30748 31297 30757 31331
rect 30757 31297 30791 31331
rect 30791 31297 30800 31331
rect 30748 31288 30800 31297
rect 31300 31288 31352 31340
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 5632 30880 5684 30932
rect 7288 30880 7340 30932
rect 8116 30923 8168 30932
rect 8116 30889 8125 30923
rect 8125 30889 8159 30923
rect 8159 30889 8168 30923
rect 8116 30880 8168 30889
rect 13544 30880 13596 30932
rect 13636 30880 13688 30932
rect 14372 30880 14424 30932
rect 16120 30880 16172 30932
rect 18788 30880 18840 30932
rect 23112 30923 23164 30932
rect 23112 30889 23121 30923
rect 23121 30889 23155 30923
rect 23155 30889 23164 30923
rect 23112 30880 23164 30889
rect 25228 30880 25280 30932
rect 8392 30812 8444 30864
rect 19156 30812 19208 30864
rect 4988 30787 5040 30796
rect 4988 30753 4997 30787
rect 4997 30753 5031 30787
rect 5031 30753 5040 30787
rect 4988 30744 5040 30753
rect 11980 30744 12032 30796
rect 12808 30744 12860 30796
rect 13544 30744 13596 30796
rect 13636 30744 13688 30796
rect 6276 30676 6328 30728
rect 7288 30719 7340 30728
rect 7288 30685 7297 30719
rect 7297 30685 7331 30719
rect 7331 30685 7340 30719
rect 7288 30676 7340 30685
rect 13268 30676 13320 30728
rect 6736 30608 6788 30660
rect 9680 30608 9732 30660
rect 14280 30608 14332 30660
rect 7932 30583 7984 30592
rect 7932 30549 7957 30583
rect 7957 30549 7984 30583
rect 7932 30540 7984 30549
rect 10232 30540 10284 30592
rect 14648 30676 14700 30728
rect 15200 30744 15252 30796
rect 17316 30787 17368 30796
rect 17316 30753 17325 30787
rect 17325 30753 17359 30787
rect 17359 30753 17368 30787
rect 17316 30744 17368 30753
rect 19524 30812 19576 30864
rect 19984 30812 20036 30864
rect 25412 30812 25464 30864
rect 22928 30744 22980 30796
rect 22284 30676 22336 30728
rect 23296 30719 23348 30728
rect 23296 30685 23305 30719
rect 23305 30685 23339 30719
rect 23339 30685 23348 30719
rect 23296 30676 23348 30685
rect 23572 30719 23624 30728
rect 23572 30685 23581 30719
rect 23581 30685 23615 30719
rect 23615 30685 23624 30719
rect 23572 30676 23624 30685
rect 26148 30744 26200 30796
rect 15200 30608 15252 30660
rect 16672 30608 16724 30660
rect 17776 30608 17828 30660
rect 19524 30608 19576 30660
rect 25044 30676 25096 30728
rect 25872 30719 25924 30728
rect 25872 30685 25881 30719
rect 25881 30685 25915 30719
rect 25915 30685 25924 30719
rect 28356 30744 28408 30796
rect 25872 30676 25924 30685
rect 28632 30676 28684 30728
rect 16212 30540 16264 30592
rect 16856 30583 16908 30592
rect 16856 30549 16865 30583
rect 16865 30549 16899 30583
rect 16899 30549 16908 30583
rect 16856 30540 16908 30549
rect 18328 30540 18380 30592
rect 19340 30540 19392 30592
rect 22284 30540 22336 30592
rect 22744 30540 22796 30592
rect 24124 30540 24176 30592
rect 24216 30540 24268 30592
rect 27712 30540 27764 30592
rect 28080 30540 28132 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 7288 30336 7340 30388
rect 12532 30336 12584 30388
rect 13452 30336 13504 30388
rect 16212 30336 16264 30388
rect 6368 30268 6420 30320
rect 6736 30268 6788 30320
rect 7932 30311 7984 30320
rect 7932 30277 7973 30311
rect 7973 30277 7984 30311
rect 7932 30268 7984 30277
rect 10876 30268 10928 30320
rect 13636 30311 13688 30320
rect 13636 30277 13645 30311
rect 13645 30277 13679 30311
rect 13679 30277 13688 30311
rect 13636 30268 13688 30277
rect 13820 30268 13872 30320
rect 14648 30268 14700 30320
rect 15200 30311 15252 30320
rect 15200 30277 15209 30311
rect 15209 30277 15243 30311
rect 15243 30277 15252 30311
rect 15200 30268 15252 30277
rect 16672 30311 16724 30320
rect 16672 30277 16681 30311
rect 16681 30277 16715 30311
rect 16715 30277 16724 30311
rect 16672 30268 16724 30277
rect 10508 30200 10560 30252
rect 15660 30200 15712 30252
rect 16948 30243 17000 30252
rect 16488 30132 16540 30184
rect 16948 30209 16957 30243
rect 16957 30209 16991 30243
rect 16991 30209 17000 30243
rect 16948 30200 17000 30209
rect 17224 30336 17276 30388
rect 17776 30379 17828 30388
rect 17776 30345 17785 30379
rect 17785 30345 17819 30379
rect 17819 30345 17828 30379
rect 17776 30336 17828 30345
rect 17132 30243 17184 30252
rect 17132 30209 17141 30243
rect 17141 30209 17175 30243
rect 17175 30209 17184 30243
rect 17132 30200 17184 30209
rect 17316 30243 17368 30252
rect 17316 30209 17325 30243
rect 17325 30209 17359 30243
rect 17359 30209 17368 30243
rect 17316 30200 17368 30209
rect 18512 30336 18564 30388
rect 18788 30379 18840 30388
rect 18788 30345 18797 30379
rect 18797 30345 18831 30379
rect 18831 30345 18840 30379
rect 18788 30336 18840 30345
rect 20812 30336 20864 30388
rect 21640 30336 21692 30388
rect 22100 30336 22152 30388
rect 23572 30336 23624 30388
rect 24952 30336 25004 30388
rect 25136 30336 25188 30388
rect 27804 30336 27856 30388
rect 28816 30336 28868 30388
rect 19340 30268 19392 30320
rect 21824 30268 21876 30320
rect 8576 30064 8628 30116
rect 12992 29996 13044 30048
rect 13636 29996 13688 30048
rect 16304 29996 16356 30048
rect 16948 29996 17000 30048
rect 18236 30243 18288 30252
rect 18236 30209 18245 30243
rect 18245 30209 18279 30243
rect 18279 30209 18288 30243
rect 18236 30200 18288 30209
rect 18512 30200 18564 30252
rect 18328 30132 18380 30184
rect 20352 30200 20404 30252
rect 24492 30268 24544 30320
rect 29184 30268 29236 30320
rect 23112 30200 23164 30252
rect 28080 30243 28132 30252
rect 28080 30209 28089 30243
rect 28089 30209 28123 30243
rect 28123 30209 28132 30243
rect 28080 30200 28132 30209
rect 22192 30132 22244 30184
rect 18328 29996 18380 30048
rect 19432 29996 19484 30048
rect 19524 29996 19576 30048
rect 25872 30064 25924 30116
rect 28080 30064 28132 30116
rect 25780 29996 25832 30048
rect 28264 29996 28316 30048
rect 28908 29996 28960 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 5816 29792 5868 29844
rect 10416 29792 10468 29844
rect 11796 29792 11848 29844
rect 12440 29792 12492 29844
rect 15752 29792 15804 29844
rect 22192 29792 22244 29844
rect 23112 29835 23164 29844
rect 23112 29801 23121 29835
rect 23121 29801 23155 29835
rect 23155 29801 23164 29835
rect 23112 29792 23164 29801
rect 24584 29792 24636 29844
rect 28908 29835 28960 29844
rect 28908 29801 28917 29835
rect 28917 29801 28951 29835
rect 28951 29801 28960 29835
rect 28908 29792 28960 29801
rect 29552 29792 29604 29844
rect 30748 29792 30800 29844
rect 9312 29656 9364 29708
rect 9772 29656 9824 29708
rect 4804 29495 4856 29504
rect 4804 29461 4813 29495
rect 4813 29461 4847 29495
rect 4847 29461 4856 29495
rect 4804 29452 4856 29461
rect 6736 29588 6788 29640
rect 8116 29588 8168 29640
rect 9036 29588 9088 29640
rect 10876 29588 10928 29640
rect 19524 29724 19576 29776
rect 22744 29724 22796 29776
rect 24768 29724 24820 29776
rect 31300 29724 31352 29776
rect 13084 29656 13136 29708
rect 13452 29656 13504 29708
rect 14924 29656 14976 29708
rect 13544 29588 13596 29640
rect 14280 29631 14332 29640
rect 5540 29520 5592 29572
rect 5908 29452 5960 29504
rect 7564 29452 7616 29504
rect 9312 29563 9364 29572
rect 9312 29529 9321 29563
rect 9321 29529 9355 29563
rect 9355 29529 9364 29563
rect 9312 29520 9364 29529
rect 10232 29520 10284 29572
rect 11612 29520 11664 29572
rect 11888 29520 11940 29572
rect 13636 29520 13688 29572
rect 14280 29597 14289 29631
rect 14289 29597 14323 29631
rect 14323 29597 14332 29631
rect 14280 29588 14332 29597
rect 14648 29588 14700 29640
rect 17316 29588 17368 29640
rect 22468 29588 22520 29640
rect 23296 29588 23348 29640
rect 24308 29656 24360 29708
rect 27528 29699 27580 29708
rect 27528 29665 27537 29699
rect 27537 29665 27571 29699
rect 27571 29665 27580 29699
rect 27528 29656 27580 29665
rect 23572 29631 23624 29640
rect 23572 29597 23581 29631
rect 23581 29597 23615 29631
rect 23615 29597 23624 29631
rect 23572 29588 23624 29597
rect 23756 29631 23808 29640
rect 23756 29597 23765 29631
rect 23765 29597 23799 29631
rect 23799 29597 23808 29631
rect 23756 29588 23808 29597
rect 24216 29588 24268 29640
rect 24676 29588 24728 29640
rect 25044 29588 25096 29640
rect 30104 29631 30156 29640
rect 30104 29597 30113 29631
rect 30113 29597 30147 29631
rect 30147 29597 30156 29631
rect 31944 29631 31996 29640
rect 30104 29588 30156 29597
rect 31944 29597 31953 29631
rect 31953 29597 31987 29631
rect 31987 29597 31996 29631
rect 31944 29588 31996 29597
rect 18512 29563 18564 29572
rect 18512 29529 18521 29563
rect 18521 29529 18555 29563
rect 18555 29529 18564 29563
rect 18512 29520 18564 29529
rect 19248 29563 19300 29572
rect 19248 29529 19257 29563
rect 19257 29529 19291 29563
rect 19291 29529 19300 29563
rect 19248 29520 19300 29529
rect 19340 29520 19392 29572
rect 20260 29520 20312 29572
rect 22744 29520 22796 29572
rect 25688 29563 25740 29572
rect 25688 29529 25722 29563
rect 25722 29529 25740 29563
rect 25688 29520 25740 29529
rect 27804 29563 27856 29572
rect 27804 29529 27838 29563
rect 27838 29529 27856 29563
rect 27804 29520 27856 29529
rect 29644 29520 29696 29572
rect 30564 29520 30616 29572
rect 10600 29452 10652 29504
rect 12072 29452 12124 29504
rect 13176 29495 13228 29504
rect 13176 29461 13185 29495
rect 13185 29461 13219 29495
rect 13219 29461 13228 29495
rect 13176 29452 13228 29461
rect 14832 29452 14884 29504
rect 21180 29452 21232 29504
rect 23756 29452 23808 29504
rect 24676 29452 24728 29504
rect 26976 29452 27028 29504
rect 30472 29452 30524 29504
rect 31300 29452 31352 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 5540 29248 5592 29300
rect 6828 29248 6880 29300
rect 10416 29291 10468 29300
rect 10416 29257 10425 29291
rect 10425 29257 10459 29291
rect 10459 29257 10468 29291
rect 10416 29248 10468 29257
rect 11612 29291 11664 29300
rect 11612 29257 11621 29291
rect 11621 29257 11655 29291
rect 11655 29257 11664 29291
rect 11612 29248 11664 29257
rect 11888 29248 11940 29300
rect 13084 29248 13136 29300
rect 14096 29291 14148 29300
rect 14096 29257 14105 29291
rect 14105 29257 14139 29291
rect 14139 29257 14148 29291
rect 14096 29248 14148 29257
rect 15844 29248 15896 29300
rect 22008 29248 22060 29300
rect 22836 29248 22888 29300
rect 23572 29248 23624 29300
rect 24584 29248 24636 29300
rect 4804 29180 4856 29232
rect 6368 29223 6420 29232
rect 6368 29189 6377 29223
rect 6377 29189 6411 29223
rect 6411 29189 6420 29223
rect 6368 29180 6420 29189
rect 6552 29223 6604 29232
rect 6552 29189 6577 29223
rect 6577 29189 6604 29223
rect 6552 29180 6604 29189
rect 7932 29180 7984 29232
rect 9036 29155 9088 29164
rect 9036 29121 9045 29155
rect 9045 29121 9079 29155
rect 9079 29121 9088 29155
rect 9036 29112 9088 29121
rect 10140 29180 10192 29232
rect 10508 29180 10560 29232
rect 10416 29112 10468 29164
rect 11796 29112 11848 29164
rect 12348 29180 12400 29232
rect 12440 29180 12492 29232
rect 12072 29155 12124 29164
rect 12072 29121 12081 29155
rect 12081 29121 12115 29155
rect 12115 29121 12124 29155
rect 12072 29112 12124 29121
rect 5816 29019 5868 29028
rect 5816 28985 5825 29019
rect 5825 28985 5859 29019
rect 5859 28985 5868 29019
rect 5816 28976 5868 28985
rect 6736 29019 6788 29028
rect 6736 28985 6745 29019
rect 6745 28985 6779 29019
rect 6779 28985 6788 29019
rect 6736 28976 6788 28985
rect 6552 28951 6604 28960
rect 6552 28917 6561 28951
rect 6561 28917 6595 28951
rect 6595 28917 6604 28951
rect 6552 28908 6604 28917
rect 11888 28908 11940 28960
rect 12808 29112 12860 29164
rect 15476 29180 15528 29232
rect 15752 29180 15804 29232
rect 14648 29112 14700 29164
rect 17776 29112 17828 29164
rect 20720 29180 20772 29232
rect 20812 29112 20864 29164
rect 21916 29180 21968 29232
rect 22192 29180 22244 29232
rect 24308 29180 24360 29232
rect 22100 29155 22152 29164
rect 22100 29121 22134 29155
rect 22134 29121 22152 29155
rect 22100 29112 22152 29121
rect 22468 29112 22520 29164
rect 23848 29155 23900 29164
rect 17408 29044 17460 29096
rect 17592 29044 17644 29096
rect 23848 29121 23857 29155
rect 23857 29121 23891 29155
rect 23891 29121 23900 29155
rect 23848 29112 23900 29121
rect 24492 29112 24544 29164
rect 24676 29112 24728 29164
rect 25688 29248 25740 29300
rect 27712 29291 27764 29300
rect 27712 29257 27721 29291
rect 27721 29257 27755 29291
rect 27755 29257 27764 29291
rect 27712 29248 27764 29257
rect 29644 29291 29696 29300
rect 29644 29257 29653 29291
rect 29653 29257 29687 29291
rect 29687 29257 29696 29291
rect 29644 29248 29696 29257
rect 30472 29248 30524 29300
rect 25780 29155 25832 29164
rect 25780 29121 25789 29155
rect 25789 29121 25823 29155
rect 25823 29121 25832 29155
rect 25780 29112 25832 29121
rect 25872 29155 25924 29164
rect 25872 29121 25881 29155
rect 25881 29121 25915 29155
rect 25915 29121 25924 29155
rect 26056 29155 26108 29164
rect 25872 29112 25924 29121
rect 26056 29121 26065 29155
rect 26065 29121 26099 29155
rect 26099 29121 26108 29155
rect 26056 29112 26108 29121
rect 29644 29112 29696 29164
rect 18512 28976 18564 29028
rect 14188 28908 14240 28960
rect 15200 28908 15252 28960
rect 15476 28908 15528 28960
rect 20536 28976 20588 29028
rect 21548 28976 21600 29028
rect 23296 28976 23348 29028
rect 25780 28976 25832 29028
rect 25964 28976 26016 29028
rect 28356 29044 28408 29096
rect 30288 29155 30340 29164
rect 29828 29044 29880 29096
rect 30288 29121 30297 29155
rect 30297 29121 30331 29155
rect 30331 29121 30340 29155
rect 30288 29112 30340 29121
rect 31024 29044 31076 29096
rect 28908 28976 28960 29028
rect 30196 28976 30248 29028
rect 30288 28976 30340 29028
rect 19892 28908 19944 28960
rect 22468 28908 22520 28960
rect 27528 28908 27580 28960
rect 27896 28908 27948 28960
rect 29920 28908 29972 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 6828 28747 6880 28756
rect 6828 28713 6837 28747
rect 6837 28713 6871 28747
rect 6871 28713 6880 28747
rect 6828 28704 6880 28713
rect 8668 28704 8720 28756
rect 12808 28704 12860 28756
rect 14648 28704 14700 28756
rect 8116 28679 8168 28688
rect 8116 28645 8125 28679
rect 8125 28645 8159 28679
rect 8159 28645 8168 28679
rect 8116 28636 8168 28645
rect 9496 28500 9548 28552
rect 14096 28568 14148 28620
rect 15016 28704 15068 28756
rect 14832 28636 14884 28688
rect 16120 28704 16172 28756
rect 20444 28704 20496 28756
rect 20812 28704 20864 28756
rect 22100 28704 22152 28756
rect 7748 28475 7800 28484
rect 7748 28441 7757 28475
rect 7757 28441 7791 28475
rect 7791 28441 7800 28475
rect 7748 28432 7800 28441
rect 7932 28475 7984 28484
rect 7932 28441 7957 28475
rect 7957 28441 7984 28475
rect 7932 28432 7984 28441
rect 12716 28432 12768 28484
rect 13176 28543 13228 28552
rect 13176 28509 13185 28543
rect 13185 28509 13219 28543
rect 13219 28509 13228 28543
rect 13176 28500 13228 28509
rect 14188 28500 14240 28552
rect 15476 28568 15528 28620
rect 15844 28500 15896 28552
rect 15476 28432 15528 28484
rect 9036 28364 9088 28416
rect 11520 28364 11572 28416
rect 12164 28364 12216 28416
rect 16764 28364 16816 28416
rect 18052 28636 18104 28688
rect 17960 28568 18012 28620
rect 18052 28543 18104 28552
rect 18052 28509 18061 28543
rect 18061 28509 18095 28543
rect 18095 28509 18104 28543
rect 18052 28500 18104 28509
rect 19800 28568 19852 28620
rect 18236 28475 18288 28484
rect 18236 28441 18245 28475
rect 18245 28441 18279 28475
rect 18279 28441 18288 28475
rect 18236 28432 18288 28441
rect 19524 28500 19576 28552
rect 19708 28543 19760 28552
rect 19708 28509 19717 28543
rect 19717 28509 19751 28543
rect 19751 28509 19760 28543
rect 19708 28500 19760 28509
rect 19892 28543 19944 28552
rect 19892 28509 19901 28543
rect 19901 28509 19935 28543
rect 19935 28509 19944 28543
rect 19892 28500 19944 28509
rect 21548 28636 21600 28688
rect 22008 28636 22060 28688
rect 23296 28704 23348 28756
rect 20536 28500 20588 28552
rect 21180 28543 21232 28552
rect 21180 28509 21189 28543
rect 21189 28509 21223 28543
rect 21223 28509 21232 28543
rect 21180 28500 21232 28509
rect 20904 28432 20956 28484
rect 21548 28500 21600 28552
rect 25872 28704 25924 28756
rect 27804 28704 27856 28756
rect 30564 28704 30616 28756
rect 31944 28704 31996 28756
rect 27528 28636 27580 28688
rect 29920 28636 29972 28688
rect 30012 28636 30064 28688
rect 30748 28636 30800 28688
rect 29736 28568 29788 28620
rect 22468 28543 22520 28552
rect 22468 28509 22477 28543
rect 22477 28509 22511 28543
rect 22511 28509 22520 28543
rect 22468 28500 22520 28509
rect 22928 28475 22980 28484
rect 22928 28441 22937 28475
rect 22937 28441 22971 28475
rect 22971 28441 22980 28475
rect 22928 28432 22980 28441
rect 18604 28364 18656 28416
rect 19064 28364 19116 28416
rect 19432 28364 19484 28416
rect 20996 28364 21048 28416
rect 21180 28364 21232 28416
rect 21824 28364 21876 28416
rect 23296 28432 23348 28484
rect 25596 28432 25648 28484
rect 26976 28475 27028 28484
rect 26976 28441 26985 28475
rect 26985 28441 27019 28475
rect 27019 28441 27028 28475
rect 26976 28432 27028 28441
rect 27896 28500 27948 28552
rect 28080 28543 28132 28552
rect 28080 28509 28089 28543
rect 28089 28509 28123 28543
rect 28123 28509 28132 28543
rect 28080 28500 28132 28509
rect 30012 28543 30064 28552
rect 30012 28509 30021 28543
rect 30021 28509 30055 28543
rect 30055 28509 30064 28543
rect 30012 28500 30064 28509
rect 23480 28364 23532 28416
rect 24216 28364 24268 28416
rect 24492 28364 24544 28416
rect 24768 28407 24820 28416
rect 24768 28373 24777 28407
rect 24777 28373 24811 28407
rect 24811 28373 24820 28407
rect 24768 28364 24820 28373
rect 26792 28364 26844 28416
rect 27988 28407 28040 28416
rect 27988 28373 27997 28407
rect 27997 28373 28031 28407
rect 28031 28373 28040 28407
rect 27988 28364 28040 28373
rect 28356 28432 28408 28484
rect 29828 28432 29880 28484
rect 30196 28543 30248 28552
rect 30196 28509 30205 28543
rect 30205 28509 30239 28543
rect 30239 28509 30248 28543
rect 30196 28500 30248 28509
rect 29000 28364 29052 28416
rect 29920 28364 29972 28416
rect 31116 28475 31168 28484
rect 31116 28441 31125 28475
rect 31125 28441 31159 28475
rect 31159 28441 31168 28475
rect 31116 28432 31168 28441
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 6368 28160 6420 28212
rect 8668 28203 8720 28212
rect 8668 28169 8677 28203
rect 8677 28169 8711 28203
rect 8711 28169 8720 28203
rect 8668 28160 8720 28169
rect 10784 28160 10836 28212
rect 13544 28160 13596 28212
rect 15476 28203 15528 28212
rect 15476 28169 15485 28203
rect 15485 28169 15519 28203
rect 15519 28169 15528 28203
rect 15476 28160 15528 28169
rect 18052 28160 18104 28212
rect 19064 28203 19116 28212
rect 19064 28169 19073 28203
rect 19073 28169 19107 28203
rect 19107 28169 19116 28203
rect 19064 28160 19116 28169
rect 20904 28160 20956 28212
rect 26332 28160 26384 28212
rect 29000 28160 29052 28212
rect 31024 28203 31076 28212
rect 7196 28024 7248 28076
rect 7564 28067 7616 28076
rect 7564 28033 7598 28067
rect 7598 28033 7616 28067
rect 7564 28024 7616 28033
rect 9036 28024 9088 28076
rect 9220 28024 9272 28076
rect 11520 28067 11572 28076
rect 11520 28033 11529 28067
rect 11529 28033 11563 28067
rect 11563 28033 11572 28067
rect 11520 28024 11572 28033
rect 11612 28024 11664 28076
rect 14924 28024 14976 28076
rect 16764 28092 16816 28144
rect 15016 27956 15068 28008
rect 16120 28067 16172 28076
rect 16120 28033 16129 28067
rect 16129 28033 16163 28067
rect 16163 28033 16172 28067
rect 16120 28024 16172 28033
rect 17500 28024 17552 28076
rect 19432 28092 19484 28144
rect 19984 28092 20036 28144
rect 24216 28135 24268 28144
rect 24216 28101 24225 28135
rect 24225 28101 24259 28135
rect 24259 28101 24268 28135
rect 24216 28092 24268 28101
rect 30380 28092 30432 28144
rect 18604 28024 18656 28076
rect 16304 27956 16356 28008
rect 17868 27956 17920 28008
rect 20260 28024 20312 28076
rect 20996 28067 21048 28076
rect 20996 28033 21005 28067
rect 21005 28033 21039 28067
rect 21039 28033 21048 28067
rect 20996 28024 21048 28033
rect 21916 28067 21968 28076
rect 21916 28033 21925 28067
rect 21925 28033 21959 28067
rect 21959 28033 21968 28067
rect 21916 28024 21968 28033
rect 22192 28067 22244 28076
rect 22192 28033 22226 28067
rect 22226 28033 22244 28067
rect 25044 28067 25096 28076
rect 22192 28024 22244 28033
rect 25044 28033 25053 28067
rect 25053 28033 25087 28067
rect 25087 28033 25096 28067
rect 25044 28024 25096 28033
rect 25320 28067 25372 28076
rect 25320 28033 25354 28067
rect 25354 28033 25372 28067
rect 25320 28024 25372 28033
rect 26976 28024 27028 28076
rect 28356 28024 28408 28076
rect 29644 28024 29696 28076
rect 29920 28067 29972 28076
rect 29920 28033 29929 28067
rect 29929 28033 29963 28067
rect 29963 28033 29972 28067
rect 29920 28024 29972 28033
rect 30196 28067 30248 28076
rect 21548 27956 21600 28008
rect 29000 27956 29052 28008
rect 30196 28033 30205 28067
rect 30205 28033 30239 28067
rect 30239 28033 30248 28067
rect 30196 28024 30248 28033
rect 31024 28169 31033 28203
rect 31033 28169 31067 28203
rect 31067 28169 31076 28203
rect 31024 28160 31076 28169
rect 31116 28092 31168 28144
rect 12716 27888 12768 27940
rect 16672 27888 16724 27940
rect 19248 27888 19300 27940
rect 19892 27888 19944 27940
rect 10508 27863 10560 27872
rect 10508 27829 10517 27863
rect 10517 27829 10551 27863
rect 10551 27829 10560 27863
rect 10508 27820 10560 27829
rect 14372 27820 14424 27872
rect 19340 27820 19392 27872
rect 19524 27820 19576 27872
rect 20168 27820 20220 27872
rect 20444 27820 20496 27872
rect 20628 27820 20680 27872
rect 20904 27820 20956 27872
rect 23388 27888 23440 27940
rect 23848 27931 23900 27940
rect 23848 27897 23857 27931
rect 23857 27897 23891 27931
rect 23891 27897 23900 27931
rect 23848 27888 23900 27897
rect 24768 27888 24820 27940
rect 29460 27888 29512 27940
rect 24308 27820 24360 27872
rect 27620 27820 27672 27872
rect 30288 27820 30340 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 6552 27616 6604 27668
rect 10508 27616 10560 27668
rect 11612 27616 11664 27668
rect 17500 27659 17552 27668
rect 10876 27548 10928 27600
rect 5448 27412 5500 27464
rect 5908 27412 5960 27464
rect 9956 27412 10008 27464
rect 10784 27412 10836 27464
rect 11428 27412 11480 27464
rect 14280 27548 14332 27600
rect 17500 27625 17509 27659
rect 17509 27625 17543 27659
rect 17543 27625 17552 27659
rect 17500 27616 17552 27625
rect 16764 27591 16816 27600
rect 11888 27455 11940 27464
rect 7748 27387 7800 27396
rect 7748 27353 7757 27387
rect 7757 27353 7791 27387
rect 7791 27353 7800 27387
rect 7748 27344 7800 27353
rect 7932 27387 7984 27396
rect 7932 27353 7957 27387
rect 7957 27353 7984 27387
rect 7932 27344 7984 27353
rect 9864 27344 9916 27396
rect 11888 27421 11897 27455
rect 11897 27421 11931 27455
rect 11931 27421 11940 27455
rect 11888 27412 11940 27421
rect 12716 27412 12768 27464
rect 14648 27480 14700 27532
rect 16764 27557 16773 27591
rect 16773 27557 16807 27591
rect 16807 27557 16816 27591
rect 16764 27548 16816 27557
rect 17408 27548 17460 27600
rect 19064 27616 19116 27668
rect 19892 27616 19944 27668
rect 20996 27616 21048 27668
rect 24032 27616 24084 27668
rect 26792 27616 26844 27668
rect 30196 27616 30248 27668
rect 13176 27344 13228 27396
rect 8116 27319 8168 27328
rect 8116 27285 8125 27319
rect 8125 27285 8159 27319
rect 8159 27285 8168 27319
rect 8116 27276 8168 27285
rect 9312 27276 9364 27328
rect 14096 27412 14148 27464
rect 19340 27548 19392 27600
rect 19708 27548 19760 27600
rect 22192 27548 22244 27600
rect 14372 27344 14424 27396
rect 14832 27344 14884 27396
rect 15292 27344 15344 27396
rect 15476 27344 15528 27396
rect 19524 27455 19576 27464
rect 19524 27421 19533 27455
rect 19533 27421 19567 27455
rect 19567 27421 19576 27455
rect 19524 27412 19576 27421
rect 18972 27344 19024 27396
rect 19708 27455 19760 27464
rect 19708 27421 19717 27455
rect 19717 27421 19751 27455
rect 19751 27421 19760 27455
rect 19708 27412 19760 27421
rect 20260 27412 20312 27464
rect 20904 27455 20956 27464
rect 20904 27421 20913 27455
rect 20913 27421 20947 27455
rect 20947 27421 20956 27455
rect 20904 27412 20956 27421
rect 21272 27412 21324 27464
rect 21364 27412 21416 27464
rect 21824 27455 21876 27464
rect 21824 27421 21833 27455
rect 21833 27421 21867 27455
rect 21867 27421 21876 27455
rect 21824 27412 21876 27421
rect 13544 27276 13596 27328
rect 13820 27276 13872 27328
rect 15844 27276 15896 27328
rect 19248 27319 19300 27328
rect 19248 27285 19257 27319
rect 19257 27285 19291 27319
rect 19291 27285 19300 27319
rect 19248 27276 19300 27285
rect 22284 27412 22336 27464
rect 23296 27548 23348 27600
rect 23848 27548 23900 27600
rect 27528 27548 27580 27600
rect 27896 27548 27948 27600
rect 28264 27548 28316 27600
rect 23204 27480 23256 27532
rect 23020 27412 23072 27464
rect 23296 27344 23348 27396
rect 24032 27344 24084 27396
rect 22284 27276 22336 27328
rect 23480 27276 23532 27328
rect 23572 27276 23624 27328
rect 24400 27387 24452 27396
rect 24400 27353 24409 27387
rect 24409 27353 24443 27387
rect 24443 27353 24452 27387
rect 24400 27344 24452 27353
rect 25872 27455 25924 27464
rect 25872 27421 25882 27455
rect 25882 27421 25916 27455
rect 25916 27421 25924 27455
rect 26148 27455 26200 27464
rect 25872 27412 25924 27421
rect 26148 27421 26157 27455
rect 26157 27421 26191 27455
rect 26191 27421 26200 27455
rect 26148 27412 26200 27421
rect 26240 27455 26292 27464
rect 26240 27421 26254 27455
rect 26254 27421 26288 27455
rect 26288 27421 26292 27455
rect 26240 27412 26292 27421
rect 26424 27412 26476 27464
rect 27804 27455 27856 27464
rect 27804 27421 27813 27455
rect 27813 27421 27847 27455
rect 27847 27421 27856 27455
rect 27804 27412 27856 27421
rect 28540 27480 28592 27532
rect 28264 27455 28316 27464
rect 28264 27421 28278 27455
rect 28278 27421 28312 27455
rect 28312 27421 28316 27455
rect 28264 27412 28316 27421
rect 26516 27344 26568 27396
rect 27712 27344 27764 27396
rect 28080 27387 28132 27396
rect 28080 27353 28089 27387
rect 28089 27353 28123 27387
rect 28123 27353 28132 27387
rect 28080 27344 28132 27353
rect 28632 27344 28684 27396
rect 29920 27548 29972 27600
rect 29736 27480 29788 27532
rect 29460 27412 29512 27464
rect 30012 27455 30064 27464
rect 30012 27421 30021 27455
rect 30021 27421 30055 27455
rect 30055 27421 30064 27455
rect 30012 27412 30064 27421
rect 31392 27344 31444 27396
rect 27252 27319 27304 27328
rect 27252 27285 27261 27319
rect 27261 27285 27295 27319
rect 27295 27285 27304 27319
rect 27252 27276 27304 27285
rect 28540 27276 28592 27328
rect 29552 27319 29604 27328
rect 29552 27285 29561 27319
rect 29561 27285 29595 27319
rect 29595 27285 29604 27319
rect 29552 27276 29604 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 5540 27004 5592 27056
rect 6920 27072 6972 27124
rect 7748 27072 7800 27124
rect 9220 27072 9272 27124
rect 10416 27115 10468 27124
rect 10416 27081 10425 27115
rect 10425 27081 10459 27115
rect 10459 27081 10468 27115
rect 10416 27072 10468 27081
rect 14280 27072 14332 27124
rect 15292 27072 15344 27124
rect 15476 27072 15528 27124
rect 6460 27004 6512 27056
rect 5448 26936 5500 26988
rect 7196 26936 7248 26988
rect 8116 26936 8168 26988
rect 8668 26979 8720 26988
rect 8668 26945 8677 26979
rect 8677 26945 8711 26979
rect 8711 26945 8720 26979
rect 8668 26936 8720 26945
rect 9956 26979 10008 26988
rect 9956 26945 9965 26979
rect 9965 26945 9999 26979
rect 9999 26945 10008 26979
rect 9956 26936 10008 26945
rect 10600 26979 10652 26988
rect 10600 26945 10609 26979
rect 10609 26945 10643 26979
rect 10643 26945 10652 26979
rect 10600 26936 10652 26945
rect 14372 26936 14424 26988
rect 14740 26936 14792 26988
rect 16764 27072 16816 27124
rect 17224 27115 17276 27124
rect 17224 27081 17233 27115
rect 17233 27081 17267 27115
rect 17267 27081 17276 27115
rect 17224 27072 17276 27081
rect 13176 26868 13228 26920
rect 13820 26868 13872 26920
rect 15108 26868 15160 26920
rect 6736 26775 6788 26784
rect 6736 26741 6745 26775
rect 6745 26741 6779 26775
rect 6779 26741 6788 26775
rect 6736 26732 6788 26741
rect 8484 26775 8536 26784
rect 8484 26741 8493 26775
rect 8493 26741 8527 26775
rect 8527 26741 8536 26775
rect 8484 26732 8536 26741
rect 9772 26775 9824 26784
rect 9772 26741 9781 26775
rect 9781 26741 9815 26775
rect 9815 26741 9824 26775
rect 9772 26732 9824 26741
rect 14280 26732 14332 26784
rect 15844 26979 15896 26988
rect 15844 26945 15853 26979
rect 15853 26945 15887 26979
rect 15887 26945 15896 26979
rect 15844 26936 15896 26945
rect 17960 26979 18012 26988
rect 17960 26945 17969 26979
rect 17969 26945 18003 26979
rect 18003 26945 18012 26979
rect 17960 26936 18012 26945
rect 19432 27004 19484 27056
rect 20628 27004 20680 27056
rect 18696 26936 18748 26988
rect 19248 26936 19300 26988
rect 19984 26936 20036 26988
rect 23848 27072 23900 27124
rect 24216 27072 24268 27124
rect 25320 27072 25372 27124
rect 23204 27047 23256 27056
rect 23204 27013 23213 27047
rect 23213 27013 23247 27047
rect 23247 27013 23256 27047
rect 23204 27004 23256 27013
rect 25872 27072 25924 27124
rect 29000 27072 29052 27124
rect 29092 27072 29144 27124
rect 20812 26868 20864 26920
rect 19984 26843 20036 26852
rect 19984 26809 19993 26843
rect 19993 26809 20027 26843
rect 20027 26809 20036 26843
rect 19984 26800 20036 26809
rect 21272 26979 21324 26988
rect 21272 26945 21281 26979
rect 21281 26945 21315 26979
rect 21315 26945 21324 26979
rect 22284 26979 22336 26988
rect 21272 26936 21324 26945
rect 22284 26945 22293 26979
rect 22293 26945 22327 26979
rect 22327 26945 22336 26979
rect 22284 26936 22336 26945
rect 22836 26936 22888 26988
rect 24032 26979 24084 26988
rect 21732 26868 21784 26920
rect 24032 26945 24041 26979
rect 24041 26945 24075 26979
rect 24075 26945 24084 26979
rect 24032 26936 24084 26945
rect 24216 26979 24268 26988
rect 24216 26945 24225 26979
rect 24225 26945 24259 26979
rect 24259 26945 24268 26979
rect 24216 26936 24268 26945
rect 25596 26936 25648 26988
rect 27252 27004 27304 27056
rect 27712 27047 27764 27056
rect 27712 27013 27721 27047
rect 27721 27013 27755 27047
rect 27755 27013 27764 27047
rect 27712 27004 27764 27013
rect 25504 26868 25556 26920
rect 22284 26800 22336 26852
rect 23296 26800 23348 26852
rect 26792 26936 26844 26988
rect 26976 26936 27028 26988
rect 27896 26979 27948 26988
rect 27896 26945 27905 26979
rect 27905 26945 27939 26979
rect 27939 26945 27948 26979
rect 28356 27004 28408 27056
rect 28908 27047 28960 27056
rect 28908 27013 28917 27047
rect 28917 27013 28951 27047
rect 28951 27013 28960 27047
rect 28908 27004 28960 27013
rect 29552 27004 29604 27056
rect 27896 26936 27948 26945
rect 26516 26868 26568 26920
rect 27804 26868 27856 26920
rect 28172 26868 28224 26920
rect 28724 26979 28776 26988
rect 28724 26945 28731 26979
rect 28731 26945 28776 26979
rect 28724 26936 28776 26945
rect 28080 26800 28132 26852
rect 16764 26732 16816 26784
rect 17776 26732 17828 26784
rect 20260 26732 20312 26784
rect 20904 26732 20956 26784
rect 23112 26732 23164 26784
rect 26240 26732 26292 26784
rect 29184 26936 29236 26988
rect 29092 26732 29144 26784
rect 30104 26732 30156 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 11520 26528 11572 26580
rect 12900 26528 12952 26580
rect 14464 26528 14516 26580
rect 13268 26460 13320 26512
rect 26240 26528 26292 26580
rect 30012 26528 30064 26580
rect 31392 26571 31444 26580
rect 31392 26537 31401 26571
rect 31401 26537 31435 26571
rect 31435 26537 31444 26571
rect 31392 26528 31444 26537
rect 5540 26324 5592 26376
rect 9036 26324 9088 26376
rect 13268 26367 13320 26376
rect 13268 26333 13277 26367
rect 13277 26333 13311 26367
rect 13311 26333 13320 26367
rect 13268 26324 13320 26333
rect 14096 26367 14148 26376
rect 5632 26256 5684 26308
rect 8484 26256 8536 26308
rect 10784 26256 10836 26308
rect 14096 26333 14105 26367
rect 14105 26333 14139 26367
rect 14139 26333 14148 26367
rect 14096 26324 14148 26333
rect 21732 26460 21784 26512
rect 24032 26460 24084 26512
rect 15200 26392 15252 26444
rect 18972 26392 19024 26444
rect 20628 26435 20680 26444
rect 20628 26401 20637 26435
rect 20637 26401 20671 26435
rect 20671 26401 20680 26435
rect 20628 26392 20680 26401
rect 23756 26392 23808 26444
rect 17960 26324 18012 26376
rect 18696 26324 18748 26376
rect 20904 26367 20956 26376
rect 20904 26333 20938 26367
rect 20938 26333 20956 26367
rect 20904 26324 20956 26333
rect 22928 26367 22980 26376
rect 22928 26333 22937 26367
rect 22937 26333 22971 26367
rect 22971 26333 22980 26367
rect 22928 26324 22980 26333
rect 6552 26188 6604 26240
rect 8392 26231 8444 26240
rect 8392 26197 8401 26231
rect 8401 26197 8435 26231
rect 8435 26197 8444 26231
rect 8392 26188 8444 26197
rect 10048 26188 10100 26240
rect 14188 26256 14240 26308
rect 15292 26256 15344 26308
rect 23112 26367 23164 26376
rect 23112 26333 23121 26367
rect 23121 26333 23155 26367
rect 23155 26333 23164 26367
rect 23112 26324 23164 26333
rect 23296 26367 23348 26376
rect 23296 26333 23305 26367
rect 23305 26333 23339 26367
rect 23339 26333 23348 26367
rect 23296 26324 23348 26333
rect 27712 26324 27764 26376
rect 29000 26324 29052 26376
rect 30104 26324 30156 26376
rect 30288 26367 30340 26376
rect 30288 26333 30322 26367
rect 30322 26333 30340 26367
rect 30288 26324 30340 26333
rect 25504 26256 25556 26308
rect 29736 26256 29788 26308
rect 14648 26188 14700 26240
rect 22744 26188 22796 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 5632 25984 5684 26036
rect 6920 25984 6972 26036
rect 6460 25916 6512 25968
rect 8668 25984 8720 26036
rect 10784 26027 10836 26036
rect 10784 25993 10793 26027
rect 10793 25993 10827 26027
rect 10827 25993 10836 26027
rect 10784 25984 10836 25993
rect 13268 25984 13320 26036
rect 14188 25984 14240 26036
rect 14464 26027 14516 26036
rect 14464 25993 14473 26027
rect 14473 25993 14507 26027
rect 14507 25993 14516 26027
rect 14464 25984 14516 25993
rect 16304 25984 16356 26036
rect 9772 25916 9824 25968
rect 16672 25916 16724 25968
rect 9036 25848 9088 25900
rect 9588 25848 9640 25900
rect 10232 25848 10284 25900
rect 13820 25848 13872 25900
rect 14280 25891 14332 25900
rect 14280 25857 14289 25891
rect 14289 25857 14323 25891
rect 14323 25857 14332 25891
rect 14280 25848 14332 25857
rect 14648 25848 14700 25900
rect 15292 25848 15344 25900
rect 16948 25984 17000 26036
rect 18420 25984 18472 26036
rect 19340 26027 19392 26036
rect 19340 25993 19349 26027
rect 19349 25993 19383 26027
rect 19383 25993 19392 26027
rect 19340 25984 19392 25993
rect 21272 25984 21324 26036
rect 24860 25984 24912 26036
rect 17316 25916 17368 25968
rect 18972 25959 19024 25968
rect 18972 25925 18981 25959
rect 18981 25925 19015 25959
rect 19015 25925 19024 25959
rect 18972 25916 19024 25925
rect 19984 25916 20036 25968
rect 17408 25848 17460 25900
rect 12532 25780 12584 25832
rect 13176 25780 13228 25832
rect 13360 25823 13412 25832
rect 13360 25789 13369 25823
rect 13369 25789 13403 25823
rect 13403 25789 13412 25823
rect 13360 25780 13412 25789
rect 14004 25780 14056 25832
rect 14188 25780 14240 25832
rect 21548 25848 21600 25900
rect 21640 25780 21692 25832
rect 25688 25848 25740 25900
rect 26240 25984 26292 26036
rect 26424 25916 26476 25968
rect 26056 25891 26108 25900
rect 26056 25857 26065 25891
rect 26065 25857 26099 25891
rect 26099 25857 26108 25891
rect 26056 25848 26108 25857
rect 25964 25780 26016 25832
rect 6552 25687 6604 25696
rect 6552 25653 6561 25687
rect 6561 25653 6595 25687
rect 6595 25653 6604 25687
rect 6552 25644 6604 25653
rect 8392 25712 8444 25764
rect 24584 25712 24636 25764
rect 26884 25848 26936 25900
rect 26424 25780 26476 25832
rect 27620 25916 27672 25968
rect 27068 25848 27120 25900
rect 29000 25916 29052 25968
rect 30472 25959 30524 25968
rect 30472 25925 30481 25959
rect 30481 25925 30515 25959
rect 30515 25925 30524 25959
rect 30472 25916 30524 25925
rect 10324 25687 10376 25696
rect 10324 25653 10333 25687
rect 10333 25653 10367 25687
rect 10367 25653 10376 25687
rect 10324 25644 10376 25653
rect 12808 25644 12860 25696
rect 17868 25644 17920 25696
rect 18788 25644 18840 25696
rect 20260 25644 20312 25696
rect 26792 25712 26844 25764
rect 30932 25848 30984 25900
rect 30380 25712 30432 25764
rect 30656 25712 30708 25764
rect 26332 25644 26384 25696
rect 28172 25644 28224 25696
rect 31024 25644 31076 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 5448 25483 5500 25492
rect 5448 25449 5457 25483
rect 5457 25449 5491 25483
rect 5491 25449 5500 25483
rect 5448 25440 5500 25449
rect 9864 25440 9916 25492
rect 10048 25483 10100 25492
rect 10048 25449 10057 25483
rect 10057 25449 10091 25483
rect 10091 25449 10100 25483
rect 10048 25440 10100 25449
rect 10232 25483 10284 25492
rect 10232 25449 10241 25483
rect 10241 25449 10275 25483
rect 10275 25449 10284 25483
rect 10232 25440 10284 25449
rect 10324 25440 10376 25492
rect 12900 25440 12952 25492
rect 17408 25483 17460 25492
rect 17408 25449 17417 25483
rect 17417 25449 17451 25483
rect 17451 25449 17460 25483
rect 17408 25440 17460 25449
rect 14924 25304 14976 25356
rect 6736 25236 6788 25288
rect 8392 25236 8444 25288
rect 9036 25236 9088 25288
rect 11980 25236 12032 25288
rect 12808 25279 12860 25288
rect 12808 25245 12817 25279
rect 12817 25245 12851 25279
rect 12851 25245 12860 25279
rect 12808 25236 12860 25245
rect 10784 25168 10836 25220
rect 17040 25236 17092 25288
rect 18420 25440 18472 25492
rect 19340 25440 19392 25492
rect 17960 25304 18012 25356
rect 19708 25304 19760 25356
rect 6644 25100 6696 25152
rect 9772 25100 9824 25152
rect 11060 25143 11112 25152
rect 11060 25109 11069 25143
rect 11069 25109 11103 25143
rect 11103 25109 11112 25143
rect 11060 25100 11112 25109
rect 11704 25100 11756 25152
rect 12164 25143 12216 25152
rect 12164 25109 12173 25143
rect 12173 25109 12207 25143
rect 12207 25109 12216 25143
rect 12164 25100 12216 25109
rect 16672 25168 16724 25220
rect 18788 25168 18840 25220
rect 19708 25168 19760 25220
rect 22008 25440 22060 25492
rect 27068 25440 27120 25492
rect 26792 25372 26844 25424
rect 30196 25372 30248 25424
rect 25964 25304 26016 25356
rect 20260 25279 20312 25288
rect 20260 25245 20269 25279
rect 20269 25245 20303 25279
rect 20303 25245 20312 25279
rect 20260 25236 20312 25245
rect 21548 25236 21600 25288
rect 22468 25279 22520 25288
rect 22468 25245 22477 25279
rect 22477 25245 22511 25279
rect 22511 25245 22520 25279
rect 22468 25236 22520 25245
rect 22744 25279 22796 25288
rect 22744 25245 22778 25279
rect 22778 25245 22796 25279
rect 22744 25236 22796 25245
rect 26424 25236 26476 25288
rect 26700 25279 26752 25288
rect 26700 25245 26709 25279
rect 26709 25245 26743 25279
rect 26743 25245 26752 25279
rect 26700 25236 26752 25245
rect 17960 25100 18012 25152
rect 24032 25168 24084 25220
rect 24860 25168 24912 25220
rect 20628 25100 20680 25152
rect 24216 25100 24268 25152
rect 24768 25100 24820 25152
rect 25780 25143 25832 25152
rect 25780 25109 25789 25143
rect 25789 25109 25823 25143
rect 25823 25109 25832 25143
rect 25780 25100 25832 25109
rect 26792 25168 26844 25220
rect 27712 25236 27764 25288
rect 27896 25279 27948 25288
rect 27896 25245 27906 25279
rect 27906 25245 27940 25279
rect 27940 25245 27948 25279
rect 28172 25279 28224 25288
rect 27896 25236 27948 25245
rect 28172 25245 28181 25279
rect 28181 25245 28215 25279
rect 28215 25245 28224 25279
rect 28172 25236 28224 25245
rect 29184 25236 29236 25288
rect 30380 25279 30432 25288
rect 30380 25245 30389 25279
rect 30389 25245 30423 25279
rect 30423 25245 30432 25279
rect 30380 25236 30432 25245
rect 31392 25304 31444 25356
rect 30748 25279 30800 25288
rect 30748 25245 30757 25279
rect 30757 25245 30791 25279
rect 30791 25245 30800 25279
rect 30748 25236 30800 25245
rect 30656 25211 30708 25220
rect 26976 25100 27028 25152
rect 30656 25177 30665 25211
rect 30665 25177 30699 25211
rect 30699 25177 30708 25211
rect 30656 25168 30708 25177
rect 28632 25100 28684 25152
rect 28908 25100 28960 25152
rect 33876 25100 33928 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 9588 24939 9640 24948
rect 9588 24905 9597 24939
rect 9597 24905 9631 24939
rect 9631 24905 9640 24939
rect 9588 24896 9640 24905
rect 12900 24939 12952 24948
rect 12900 24905 12909 24939
rect 12909 24905 12943 24939
rect 12943 24905 12952 24939
rect 12900 24896 12952 24905
rect 6920 24871 6972 24880
rect 6920 24837 6929 24871
rect 6929 24837 6963 24871
rect 6963 24837 6972 24871
rect 6920 24828 6972 24837
rect 4712 24803 4764 24812
rect 4712 24769 4721 24803
rect 4721 24769 4755 24803
rect 4755 24769 4764 24803
rect 4712 24760 4764 24769
rect 6184 24760 6236 24812
rect 11060 24828 11112 24880
rect 12164 24828 12216 24880
rect 13544 24828 13596 24880
rect 13636 24803 13688 24812
rect 13636 24769 13645 24803
rect 13645 24769 13679 24803
rect 13679 24769 13688 24803
rect 13636 24760 13688 24769
rect 4620 24556 4672 24608
rect 7104 24599 7156 24608
rect 7104 24565 7113 24599
rect 7113 24565 7147 24599
rect 7147 24565 7156 24599
rect 7104 24556 7156 24565
rect 7288 24599 7340 24608
rect 7288 24565 7297 24599
rect 7297 24565 7331 24599
rect 7331 24565 7340 24599
rect 7288 24556 7340 24565
rect 13360 24692 13412 24744
rect 13820 24803 13872 24812
rect 13820 24769 13829 24803
rect 13829 24769 13863 24803
rect 13863 24769 13872 24803
rect 16672 24828 16724 24880
rect 13820 24760 13872 24769
rect 14280 24760 14332 24812
rect 14464 24692 14516 24744
rect 16856 24760 16908 24812
rect 14004 24556 14056 24608
rect 14096 24556 14148 24608
rect 16764 24692 16816 24744
rect 17132 24803 17184 24812
rect 17132 24769 17141 24803
rect 17141 24769 17175 24803
rect 17175 24769 17184 24803
rect 17132 24760 17184 24769
rect 17776 24760 17828 24812
rect 17960 24760 18012 24812
rect 19064 24896 19116 24948
rect 20720 24896 20772 24948
rect 21180 24896 21232 24948
rect 22100 24896 22152 24948
rect 24032 24939 24084 24948
rect 19984 24871 20036 24880
rect 18972 24760 19024 24812
rect 19432 24760 19484 24812
rect 19984 24837 20018 24871
rect 20018 24837 20036 24871
rect 19984 24828 20036 24837
rect 22560 24828 22612 24880
rect 24032 24905 24041 24939
rect 24041 24905 24075 24939
rect 24075 24905 24084 24939
rect 24032 24896 24084 24905
rect 22652 24760 22704 24812
rect 17316 24624 17368 24676
rect 19340 24692 19392 24744
rect 25780 24896 25832 24948
rect 26700 24896 26752 24948
rect 27896 24896 27948 24948
rect 29184 24896 29236 24948
rect 30472 24896 30524 24948
rect 24860 24828 24912 24880
rect 26608 24828 26660 24880
rect 24492 24803 24544 24812
rect 24492 24769 24501 24803
rect 24501 24769 24535 24803
rect 24535 24769 24544 24803
rect 24676 24803 24728 24812
rect 24492 24760 24544 24769
rect 24676 24769 24685 24803
rect 24685 24769 24719 24803
rect 24719 24769 24728 24803
rect 24676 24760 24728 24769
rect 25964 24803 26016 24812
rect 23020 24692 23072 24744
rect 25964 24769 25973 24803
rect 25973 24769 26007 24803
rect 26007 24769 26016 24803
rect 25964 24760 26016 24769
rect 26792 24760 26844 24812
rect 27068 24760 27120 24812
rect 28908 24828 28960 24880
rect 30196 24828 30248 24880
rect 26424 24692 26476 24744
rect 16856 24556 16908 24608
rect 17960 24556 18012 24608
rect 18972 24556 19024 24608
rect 19524 24556 19576 24608
rect 25136 24624 25188 24676
rect 26516 24624 26568 24676
rect 26884 24624 26936 24676
rect 30564 24803 30616 24812
rect 30564 24769 30573 24803
rect 30573 24769 30607 24803
rect 30607 24769 30616 24803
rect 30564 24760 30616 24769
rect 30840 24760 30892 24812
rect 31392 24803 31444 24812
rect 30656 24692 30708 24744
rect 31392 24769 31401 24803
rect 31401 24769 31435 24803
rect 31435 24769 31444 24803
rect 31392 24760 31444 24769
rect 31208 24667 31260 24676
rect 31208 24633 31217 24667
rect 31217 24633 31251 24667
rect 31251 24633 31260 24667
rect 31208 24624 31260 24633
rect 22744 24556 22796 24608
rect 25964 24556 26016 24608
rect 29000 24556 29052 24608
rect 31116 24556 31168 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 7104 24352 7156 24404
rect 7748 24352 7800 24404
rect 8392 24395 8444 24404
rect 8392 24361 8401 24395
rect 8401 24361 8435 24395
rect 8435 24361 8444 24395
rect 8392 24352 8444 24361
rect 9588 24352 9640 24404
rect 9956 24352 10008 24404
rect 10140 24284 10192 24336
rect 13820 24284 13872 24336
rect 5540 24216 5592 24268
rect 12808 24216 12860 24268
rect 14464 24216 14516 24268
rect 4620 24080 4672 24132
rect 6736 24080 6788 24132
rect 6920 24080 6972 24132
rect 7380 24080 7432 24132
rect 11520 24148 11572 24200
rect 14648 24148 14700 24200
rect 15568 24191 15620 24200
rect 15568 24157 15577 24191
rect 15577 24157 15611 24191
rect 15611 24157 15620 24191
rect 15568 24148 15620 24157
rect 24308 24284 24360 24336
rect 24492 24352 24544 24404
rect 27068 24352 27120 24404
rect 28448 24352 28500 24404
rect 18328 24216 18380 24268
rect 19340 24216 19392 24268
rect 19524 24191 19576 24200
rect 19524 24157 19533 24191
rect 19533 24157 19567 24191
rect 19567 24157 19576 24191
rect 19524 24148 19576 24157
rect 20720 24216 20772 24268
rect 23204 24216 23256 24268
rect 19708 24191 19760 24200
rect 19708 24157 19717 24191
rect 19717 24157 19751 24191
rect 19751 24157 19760 24191
rect 19708 24148 19760 24157
rect 19984 24148 20036 24200
rect 20260 24148 20312 24200
rect 21548 24148 21600 24200
rect 22100 24148 22152 24200
rect 25964 24284 26016 24336
rect 26884 24284 26936 24336
rect 30932 24352 30984 24404
rect 31392 24352 31444 24404
rect 11796 24080 11848 24132
rect 16212 24080 16264 24132
rect 17316 24123 17368 24132
rect 17316 24089 17325 24123
rect 17325 24089 17359 24123
rect 17359 24089 17368 24123
rect 17316 24080 17368 24089
rect 20628 24123 20680 24132
rect 5356 24012 5408 24064
rect 6184 24012 6236 24064
rect 8576 24012 8628 24064
rect 9036 24012 9088 24064
rect 9312 24055 9364 24064
rect 9312 24021 9321 24055
rect 9321 24021 9355 24055
rect 9355 24021 9364 24055
rect 9312 24012 9364 24021
rect 10140 24012 10192 24064
rect 19294 24012 19346 24064
rect 20628 24089 20637 24123
rect 20637 24089 20671 24123
rect 20671 24089 20680 24123
rect 20628 24080 20680 24089
rect 21180 24123 21232 24132
rect 21180 24089 21189 24123
rect 21189 24089 21223 24123
rect 21223 24089 21232 24123
rect 21180 24080 21232 24089
rect 21640 24080 21692 24132
rect 22652 24080 22704 24132
rect 24860 24148 24912 24200
rect 25044 24148 25096 24200
rect 26792 24191 26844 24200
rect 26792 24157 26801 24191
rect 26801 24157 26835 24191
rect 26835 24157 26844 24191
rect 26792 24148 26844 24157
rect 28908 24216 28960 24268
rect 31116 24216 31168 24268
rect 25320 24080 25372 24132
rect 26148 24080 26200 24132
rect 26700 24080 26752 24132
rect 22836 24012 22888 24064
rect 23756 24055 23808 24064
rect 23756 24021 23765 24055
rect 23765 24021 23799 24055
rect 23799 24021 23808 24055
rect 23756 24012 23808 24021
rect 25688 24012 25740 24064
rect 28448 24148 28500 24200
rect 30104 24148 30156 24200
rect 28264 24080 28316 24132
rect 28356 24012 28408 24064
rect 28724 24012 28776 24064
rect 30288 24012 30340 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 4712 23808 4764 23860
rect 4896 23672 4948 23724
rect 6184 23740 6236 23792
rect 6920 23808 6972 23860
rect 7748 23851 7800 23860
rect 7748 23817 7757 23851
rect 7757 23817 7791 23851
rect 7791 23817 7800 23851
rect 7748 23808 7800 23817
rect 9588 23851 9640 23860
rect 9588 23817 9597 23851
rect 9597 23817 9631 23851
rect 9631 23817 9640 23851
rect 9588 23808 9640 23817
rect 10784 23808 10836 23860
rect 11520 23808 11572 23860
rect 17132 23808 17184 23860
rect 6644 23715 6696 23724
rect 6644 23681 6678 23715
rect 6678 23681 6696 23715
rect 6644 23672 6696 23681
rect 11704 23783 11756 23792
rect 11704 23749 11713 23783
rect 11713 23749 11747 23783
rect 11747 23749 11756 23783
rect 11704 23740 11756 23749
rect 14004 23740 14056 23792
rect 14648 23740 14700 23792
rect 17316 23740 17368 23792
rect 19524 23783 19576 23792
rect 8300 23672 8352 23724
rect 8484 23715 8536 23724
rect 8484 23681 8518 23715
rect 8518 23681 8536 23715
rect 8484 23672 8536 23681
rect 11428 23672 11480 23724
rect 13357 23718 13409 23727
rect 13357 23684 13384 23718
rect 13384 23684 13409 23718
rect 13357 23675 13409 23684
rect 13912 23672 13964 23724
rect 14096 23715 14148 23724
rect 14096 23681 14105 23715
rect 14105 23681 14139 23715
rect 14139 23681 14148 23715
rect 14096 23672 14148 23681
rect 13268 23536 13320 23588
rect 14004 23604 14056 23656
rect 16212 23536 16264 23588
rect 4620 23468 4672 23520
rect 5356 23511 5408 23520
rect 5356 23477 5365 23511
rect 5365 23477 5399 23511
rect 5399 23477 5408 23511
rect 5356 23468 5408 23477
rect 10600 23511 10652 23520
rect 10600 23477 10609 23511
rect 10609 23477 10643 23511
rect 10643 23477 10652 23511
rect 10600 23468 10652 23477
rect 10784 23511 10836 23520
rect 10784 23477 10793 23511
rect 10793 23477 10827 23511
rect 10827 23477 10836 23511
rect 10784 23468 10836 23477
rect 13084 23468 13136 23520
rect 17500 23672 17552 23724
rect 19524 23749 19536 23783
rect 19536 23749 19576 23783
rect 19524 23740 19576 23749
rect 19984 23740 20036 23792
rect 22560 23740 22612 23792
rect 22836 23808 22888 23860
rect 23296 23808 23348 23860
rect 25136 23808 25188 23860
rect 25780 23808 25832 23860
rect 26056 23808 26108 23860
rect 28264 23851 28316 23860
rect 28264 23817 28273 23851
rect 28273 23817 28307 23851
rect 28307 23817 28316 23851
rect 28264 23808 28316 23817
rect 28724 23808 28776 23860
rect 30564 23808 30616 23860
rect 22100 23715 22152 23724
rect 22100 23681 22109 23715
rect 22109 23681 22143 23715
rect 22143 23681 22152 23715
rect 22100 23672 22152 23681
rect 22652 23672 22704 23724
rect 24308 23740 24360 23792
rect 25044 23672 25096 23724
rect 25320 23715 25372 23724
rect 25320 23681 25329 23715
rect 25329 23681 25363 23715
rect 25363 23681 25372 23715
rect 25320 23672 25372 23681
rect 26700 23740 26752 23792
rect 25504 23715 25556 23724
rect 25504 23681 25513 23715
rect 25513 23681 25547 23715
rect 25547 23681 25556 23715
rect 25504 23672 25556 23681
rect 25688 23715 25740 23724
rect 25688 23681 25697 23715
rect 25697 23681 25731 23715
rect 25731 23681 25740 23715
rect 26148 23715 26200 23724
rect 25688 23672 25740 23681
rect 26148 23681 26157 23715
rect 26157 23681 26191 23715
rect 26191 23681 26200 23715
rect 26148 23672 26200 23681
rect 26424 23672 26476 23724
rect 20996 23604 21048 23656
rect 25872 23604 25924 23656
rect 27896 23672 27948 23724
rect 28080 23672 28132 23724
rect 28264 23672 28316 23724
rect 28724 23715 28776 23724
rect 28724 23681 28733 23715
rect 28733 23681 28767 23715
rect 28767 23681 28776 23715
rect 30288 23740 30340 23792
rect 28724 23672 28776 23681
rect 29000 23672 29052 23724
rect 29736 23672 29788 23724
rect 30380 23715 30432 23724
rect 30380 23681 30389 23715
rect 30389 23681 30423 23715
rect 30423 23681 30432 23715
rect 30380 23672 30432 23681
rect 31392 23740 31444 23792
rect 18880 23536 18932 23588
rect 20444 23536 20496 23588
rect 22100 23536 22152 23588
rect 22284 23536 22336 23588
rect 24400 23536 24452 23588
rect 27160 23536 27212 23588
rect 30380 23536 30432 23588
rect 18696 23468 18748 23520
rect 19156 23468 19208 23520
rect 22008 23468 22060 23520
rect 23112 23468 23164 23520
rect 27712 23468 27764 23520
rect 28448 23468 28500 23520
rect 30564 23672 30616 23724
rect 30932 23672 30984 23724
rect 30748 23604 30800 23656
rect 31668 23468 31720 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 6736 23307 6788 23316
rect 6736 23273 6745 23307
rect 6745 23273 6779 23307
rect 6779 23273 6788 23307
rect 6736 23264 6788 23273
rect 8484 23264 8536 23316
rect 10600 23264 10652 23316
rect 11704 23264 11756 23316
rect 14004 23264 14056 23316
rect 17500 23264 17552 23316
rect 18604 23307 18656 23316
rect 18604 23273 18613 23307
rect 18613 23273 18647 23307
rect 18647 23273 18656 23307
rect 18604 23264 18656 23273
rect 17224 23196 17276 23248
rect 18880 23196 18932 23248
rect 21180 23264 21232 23316
rect 25504 23264 25556 23316
rect 26240 23307 26292 23316
rect 26240 23273 26249 23307
rect 26249 23273 26283 23307
rect 26283 23273 26292 23307
rect 26240 23264 26292 23273
rect 28724 23264 28776 23316
rect 30012 23264 30064 23316
rect 30564 23264 30616 23316
rect 22192 23196 22244 23248
rect 8300 23128 8352 23180
rect 8944 23128 8996 23180
rect 3792 23103 3844 23112
rect 3792 23069 3801 23103
rect 3801 23069 3835 23103
rect 3835 23069 3844 23103
rect 3792 23060 3844 23069
rect 4620 23060 4672 23112
rect 7288 23060 7340 23112
rect 9220 23060 9272 23112
rect 11796 23060 11848 23112
rect 14648 23060 14700 23112
rect 16120 23103 16172 23112
rect 16120 23069 16129 23103
rect 16129 23069 16163 23103
rect 16163 23069 16172 23103
rect 16120 23060 16172 23069
rect 16396 23060 16448 23112
rect 17224 23060 17276 23112
rect 10048 22992 10100 23044
rect 13452 22992 13504 23044
rect 16672 22992 16724 23044
rect 18328 23060 18380 23112
rect 18604 23060 18656 23112
rect 20720 23128 20772 23180
rect 20260 23060 20312 23112
rect 20812 23060 20864 23112
rect 23756 23128 23808 23180
rect 20904 23035 20956 23044
rect 4712 22924 4764 22976
rect 12348 22924 12400 22976
rect 20260 22924 20312 22976
rect 20904 23001 20913 23035
rect 20913 23001 20947 23035
rect 20947 23001 20956 23035
rect 20904 22992 20956 23001
rect 22284 23103 22336 23112
rect 22284 23069 22293 23103
rect 22293 23069 22327 23103
rect 22327 23069 22336 23103
rect 22284 23060 22336 23069
rect 22560 23060 22612 23112
rect 23388 23060 23440 23112
rect 25044 23060 25096 23112
rect 26424 23060 26476 23112
rect 28448 23060 28500 23112
rect 32680 23103 32732 23112
rect 32680 23069 32689 23103
rect 32689 23069 32723 23103
rect 32723 23069 32732 23103
rect 32680 23060 32732 23069
rect 23480 22992 23532 23044
rect 25780 22992 25832 23044
rect 21180 22924 21232 22976
rect 21916 22924 21968 22976
rect 22192 22924 22244 22976
rect 22560 22924 22612 22976
rect 32496 22967 32548 22976
rect 32496 22933 32505 22967
rect 32505 22933 32539 22967
rect 32539 22933 32548 22967
rect 32496 22924 32548 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 20 22516 72 22568
rect 5448 22652 5500 22704
rect 5724 22584 5776 22636
rect 7840 22652 7892 22704
rect 11520 22695 11572 22704
rect 11520 22661 11529 22695
rect 11529 22661 11563 22695
rect 11563 22661 11572 22695
rect 11520 22652 11572 22661
rect 11704 22695 11756 22704
rect 11704 22661 11729 22695
rect 11729 22661 11756 22695
rect 13452 22720 13504 22772
rect 18144 22720 18196 22772
rect 19984 22720 20036 22772
rect 23480 22720 23532 22772
rect 23940 22720 23992 22772
rect 26424 22763 26476 22772
rect 26424 22729 26433 22763
rect 26433 22729 26467 22763
rect 26467 22729 26476 22763
rect 26424 22720 26476 22729
rect 11704 22652 11756 22661
rect 7196 22584 7248 22636
rect 8668 22584 8720 22636
rect 10784 22584 10836 22636
rect 11244 22584 11296 22636
rect 12900 22584 12952 22636
rect 13084 22584 13136 22636
rect 18236 22584 18288 22636
rect 19248 22584 19300 22636
rect 22468 22652 22520 22704
rect 21916 22584 21968 22636
rect 23480 22584 23532 22636
rect 23848 22627 23900 22636
rect 8576 22559 8628 22568
rect 8576 22525 8585 22559
rect 8585 22525 8619 22559
rect 8619 22525 8628 22559
rect 8576 22516 8628 22525
rect 12440 22516 12492 22568
rect 18788 22516 18840 22568
rect 23848 22593 23857 22627
rect 23857 22593 23891 22627
rect 23891 22593 23900 22627
rect 23848 22584 23900 22593
rect 25044 22627 25096 22636
rect 25044 22593 25053 22627
rect 25053 22593 25087 22627
rect 25087 22593 25096 22627
rect 25044 22584 25096 22593
rect 25136 22584 25188 22636
rect 29276 22652 29328 22704
rect 23756 22516 23808 22568
rect 27344 22516 27396 22568
rect 27896 22627 27948 22636
rect 27896 22593 27905 22627
rect 27905 22593 27939 22627
rect 27939 22593 27948 22627
rect 27896 22584 27948 22593
rect 28356 22584 28408 22636
rect 29920 22584 29972 22636
rect 30564 22652 30616 22704
rect 30932 22584 30984 22636
rect 32496 22652 32548 22704
rect 34152 22627 34204 22636
rect 34152 22593 34161 22627
rect 34161 22593 34195 22627
rect 34195 22593 34204 22627
rect 34152 22584 34204 22593
rect 4896 22491 4948 22500
rect 4896 22457 4905 22491
rect 4905 22457 4939 22491
rect 4939 22457 4948 22491
rect 4896 22448 4948 22457
rect 4712 22423 4764 22432
rect 4712 22389 4721 22423
rect 4721 22389 4755 22423
rect 4755 22389 4764 22423
rect 4712 22380 4764 22389
rect 7012 22448 7064 22500
rect 7380 22491 7432 22500
rect 7380 22457 7389 22491
rect 7389 22457 7423 22491
rect 7423 22457 7432 22491
rect 7380 22448 7432 22457
rect 10048 22491 10100 22500
rect 10048 22457 10057 22491
rect 10057 22457 10091 22491
rect 10091 22457 10100 22491
rect 10048 22448 10100 22457
rect 6920 22423 6972 22432
rect 6920 22389 6929 22423
rect 6929 22389 6963 22423
rect 6963 22389 6972 22423
rect 6920 22380 6972 22389
rect 12164 22448 12216 22500
rect 17776 22448 17828 22500
rect 20720 22448 20772 22500
rect 11888 22423 11940 22432
rect 11888 22389 11897 22423
rect 11897 22389 11931 22423
rect 11931 22389 11940 22423
rect 11888 22380 11940 22389
rect 12348 22423 12400 22432
rect 12348 22389 12357 22423
rect 12357 22389 12391 22423
rect 12391 22389 12400 22423
rect 12348 22380 12400 22389
rect 17500 22380 17552 22432
rect 18144 22380 18196 22432
rect 27712 22380 27764 22432
rect 28080 22380 28132 22432
rect 28908 22380 28960 22432
rect 31300 22380 31352 22432
rect 33508 22423 33560 22432
rect 33508 22389 33517 22423
rect 33517 22389 33551 22423
rect 33551 22389 33560 22423
rect 33508 22380 33560 22389
rect 33968 22423 34020 22432
rect 33968 22389 33977 22423
rect 33977 22389 34011 22423
rect 34011 22389 34020 22423
rect 33968 22380 34020 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 7012 22219 7064 22228
rect 7012 22185 7021 22219
rect 7021 22185 7055 22219
rect 7055 22185 7064 22219
rect 7012 22176 7064 22185
rect 8668 22176 8720 22228
rect 12164 22219 12216 22228
rect 12164 22185 12173 22219
rect 12173 22185 12207 22219
rect 12207 22185 12216 22219
rect 12164 22176 12216 22185
rect 12808 22219 12860 22228
rect 12808 22185 12817 22219
rect 12817 22185 12851 22219
rect 12851 22185 12860 22219
rect 12808 22176 12860 22185
rect 12900 22176 12952 22228
rect 13084 22176 13136 22228
rect 18236 22176 18288 22228
rect 19156 22176 19208 22228
rect 20904 22176 20956 22228
rect 21548 22176 21600 22228
rect 20812 22108 20864 22160
rect 5448 22040 5500 22092
rect 3792 21972 3844 22024
rect 8668 22040 8720 22092
rect 12900 22040 12952 22092
rect 10876 21972 10928 22024
rect 12440 21972 12492 22024
rect 14096 21972 14148 22024
rect 17960 22040 18012 22092
rect 22468 22083 22520 22092
rect 15660 21972 15712 22024
rect 17316 21972 17368 22024
rect 22468 22049 22477 22083
rect 22477 22049 22511 22083
rect 22511 22049 22520 22083
rect 22468 22040 22520 22049
rect 23940 22040 23992 22092
rect 6276 21904 6328 21956
rect 11336 21904 11388 21956
rect 11520 21904 11572 21956
rect 15568 21904 15620 21956
rect 16212 21904 16264 21956
rect 19064 21904 19116 21956
rect 20076 21947 20128 21956
rect 20076 21913 20110 21947
rect 20110 21913 20128 21947
rect 20076 21904 20128 21913
rect 22100 21904 22152 21956
rect 22836 21904 22888 21956
rect 24768 22015 24820 22024
rect 24768 21981 24775 22015
rect 24775 21981 24820 22015
rect 24768 21972 24820 21981
rect 24952 22015 25004 22024
rect 24952 21981 24961 22015
rect 24961 21981 24995 22015
rect 24995 21981 25004 22015
rect 24952 21972 25004 21981
rect 25136 21972 25188 22024
rect 25780 22108 25832 22160
rect 26424 22108 26476 22160
rect 26516 22040 26568 22092
rect 28448 22176 28500 22228
rect 28908 22176 28960 22228
rect 30932 22219 30984 22228
rect 30932 22185 30941 22219
rect 30941 22185 30975 22219
rect 30975 22185 30984 22219
rect 30932 22176 30984 22185
rect 30104 22108 30156 22160
rect 30196 22108 30248 22160
rect 29828 22083 29880 22092
rect 29828 22049 29837 22083
rect 29837 22049 29871 22083
rect 29871 22049 29880 22083
rect 29828 22040 29880 22049
rect 26056 22015 26108 22024
rect 26056 21981 26065 22015
rect 26065 21981 26099 22015
rect 26099 21981 26108 22015
rect 26056 21972 26108 21981
rect 26148 22015 26200 22024
rect 26148 21981 26162 22015
rect 26162 21981 26196 22015
rect 26196 21981 26200 22015
rect 26148 21972 26200 21981
rect 26608 21972 26660 22024
rect 27692 21947 27744 21956
rect 27692 21913 27701 21947
rect 27701 21913 27735 21947
rect 27735 21913 27744 21947
rect 28816 21972 28868 22024
rect 30748 22040 30800 22092
rect 27692 21904 27744 21913
rect 29920 21904 29972 21956
rect 30472 22015 30524 22024
rect 30472 21981 30481 22015
rect 30481 21981 30515 22015
rect 30515 21981 30524 22015
rect 30472 21972 30524 21981
rect 30840 21972 30892 22024
rect 31208 22015 31260 22024
rect 31208 21981 31217 22015
rect 31217 21981 31251 22015
rect 31251 21981 31260 22015
rect 31208 21972 31260 21981
rect 30656 21904 30708 21956
rect 31392 22015 31444 22024
rect 31392 21981 31401 22015
rect 31401 21981 31435 22015
rect 31435 21981 31444 22015
rect 33508 22040 33560 22092
rect 31392 21972 31444 21981
rect 31668 21972 31720 22024
rect 32864 22015 32916 22024
rect 32864 21981 32873 22015
rect 32873 21981 32907 22015
rect 32907 21981 32916 22015
rect 32864 21972 32916 21981
rect 34980 21972 35032 22024
rect 11244 21836 11296 21888
rect 13084 21836 13136 21888
rect 15200 21836 15252 21888
rect 16304 21836 16356 21888
rect 16856 21836 16908 21888
rect 17960 21836 18012 21888
rect 18696 21879 18748 21888
rect 18696 21845 18705 21879
rect 18705 21845 18739 21879
rect 18739 21845 18748 21879
rect 18696 21836 18748 21845
rect 21732 21836 21784 21888
rect 23848 21879 23900 21888
rect 23848 21845 23857 21879
rect 23857 21845 23891 21879
rect 23891 21845 23900 21879
rect 23848 21836 23900 21845
rect 24584 21836 24636 21888
rect 25320 21836 25372 21888
rect 25780 21836 25832 21888
rect 32772 21836 32824 21888
rect 33784 21836 33836 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 7564 21632 7616 21684
rect 7840 21675 7892 21684
rect 7840 21641 7865 21675
rect 7865 21641 7892 21675
rect 7840 21632 7892 21641
rect 12808 21632 12860 21684
rect 15568 21675 15620 21684
rect 15568 21641 15577 21675
rect 15577 21641 15611 21675
rect 15611 21641 15620 21675
rect 15568 21632 15620 21641
rect 15660 21632 15712 21684
rect 18604 21632 18656 21684
rect 18788 21675 18840 21684
rect 18788 21641 18797 21675
rect 18797 21641 18831 21675
rect 18831 21641 18840 21675
rect 18788 21632 18840 21641
rect 19064 21632 19116 21684
rect 7380 21564 7432 21616
rect 12348 21564 12400 21616
rect 5080 21539 5132 21548
rect 5080 21505 5089 21539
rect 5089 21505 5123 21539
rect 5123 21505 5132 21539
rect 5080 21496 5132 21505
rect 7012 21496 7064 21548
rect 8668 21539 8720 21548
rect 8668 21505 8677 21539
rect 8677 21505 8711 21539
rect 8711 21505 8720 21539
rect 8668 21496 8720 21505
rect 9220 21539 9272 21548
rect 9220 21505 9229 21539
rect 9229 21505 9263 21539
rect 9263 21505 9272 21539
rect 9220 21496 9272 21505
rect 14924 21539 14976 21548
rect 14924 21505 14933 21539
rect 14933 21505 14967 21539
rect 14967 21505 14976 21539
rect 14924 21496 14976 21505
rect 15752 21539 15804 21548
rect 15752 21505 15761 21539
rect 15761 21505 15795 21539
rect 15795 21505 15804 21539
rect 15752 21496 15804 21505
rect 15844 21539 15896 21548
rect 15844 21505 15853 21539
rect 15853 21505 15887 21539
rect 15887 21505 15896 21539
rect 16488 21564 16540 21616
rect 19248 21564 19300 21616
rect 22652 21632 22704 21684
rect 22836 21675 22888 21684
rect 22836 21641 22845 21675
rect 22845 21641 22879 21675
rect 22879 21641 22888 21675
rect 22836 21632 22888 21641
rect 23112 21632 23164 21684
rect 22744 21564 22796 21616
rect 25044 21632 25096 21684
rect 27712 21632 27764 21684
rect 15844 21496 15896 21505
rect 5724 21428 5776 21480
rect 6460 21428 6512 21480
rect 10876 21428 10928 21480
rect 15200 21428 15252 21480
rect 17316 21496 17368 21548
rect 18420 21496 18472 21548
rect 18696 21496 18748 21548
rect 23664 21564 23716 21616
rect 28264 21632 28316 21684
rect 29920 21632 29972 21684
rect 28448 21564 28500 21616
rect 29552 21564 29604 21616
rect 4620 21292 4672 21344
rect 4896 21335 4948 21344
rect 4896 21301 4905 21335
rect 4905 21301 4939 21335
rect 4939 21301 4948 21335
rect 4896 21292 4948 21301
rect 9496 21360 9548 21412
rect 15568 21360 15620 21412
rect 16764 21428 16816 21480
rect 17132 21428 17184 21480
rect 20904 21428 20956 21480
rect 23388 21496 23440 21548
rect 24032 21539 24084 21548
rect 24032 21505 24041 21539
rect 24041 21505 24075 21539
rect 24075 21505 24084 21539
rect 24032 21496 24084 21505
rect 27160 21496 27212 21548
rect 23664 21428 23716 21480
rect 27436 21496 27488 21548
rect 27896 21539 27948 21548
rect 27896 21505 27905 21539
rect 27905 21505 27939 21539
rect 27939 21505 27948 21539
rect 27896 21496 27948 21505
rect 24584 21360 24636 21412
rect 28080 21360 28132 21412
rect 28356 21539 28408 21548
rect 28356 21505 28370 21539
rect 28370 21505 28404 21539
rect 28404 21505 28408 21539
rect 29000 21539 29052 21548
rect 28356 21496 28408 21505
rect 29000 21505 29009 21539
rect 29009 21505 29043 21539
rect 29043 21505 29052 21539
rect 29000 21496 29052 21505
rect 29276 21496 29328 21548
rect 29736 21496 29788 21548
rect 30104 21632 30156 21684
rect 31576 21632 31628 21684
rect 32680 21675 32732 21684
rect 32680 21641 32689 21675
rect 32689 21641 32723 21675
rect 32723 21641 32732 21675
rect 32680 21632 32732 21641
rect 34980 21675 35032 21684
rect 34980 21641 34989 21675
rect 34989 21641 35023 21675
rect 35023 21641 35032 21675
rect 34980 21632 35032 21641
rect 30104 21539 30156 21548
rect 30104 21505 30113 21539
rect 30113 21505 30147 21539
rect 30147 21505 30156 21539
rect 30104 21496 30156 21505
rect 30472 21496 30524 21548
rect 30932 21539 30984 21548
rect 30932 21505 30941 21539
rect 30941 21505 30975 21539
rect 30975 21505 30984 21539
rect 30932 21496 30984 21505
rect 33508 21564 33560 21616
rect 33968 21564 34020 21616
rect 31944 21496 31996 21548
rect 32772 21496 32824 21548
rect 31392 21428 31444 21480
rect 33600 21471 33652 21480
rect 33600 21437 33609 21471
rect 33609 21437 33643 21471
rect 33643 21437 33652 21471
rect 33600 21428 33652 21437
rect 31208 21360 31260 21412
rect 8300 21292 8352 21344
rect 8944 21292 8996 21344
rect 22100 21335 22152 21344
rect 22100 21301 22109 21335
rect 22109 21301 22143 21335
rect 22143 21301 22152 21335
rect 22100 21292 22152 21301
rect 24400 21292 24452 21344
rect 25596 21292 25648 21344
rect 27068 21292 27120 21344
rect 28264 21292 28316 21344
rect 30472 21335 30524 21344
rect 30472 21301 30481 21335
rect 30481 21301 30515 21335
rect 30515 21301 30524 21335
rect 30472 21292 30524 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 6276 21131 6328 21140
rect 6276 21097 6285 21131
rect 6285 21097 6319 21131
rect 6319 21097 6328 21131
rect 6276 21088 6328 21097
rect 3792 20927 3844 20936
rect 3792 20893 3801 20927
rect 3801 20893 3835 20927
rect 3835 20893 3844 20927
rect 3792 20884 3844 20893
rect 4896 20884 4948 20936
rect 6920 20884 6972 20936
rect 7380 20859 7432 20868
rect 7380 20825 7389 20859
rect 7389 20825 7423 20859
rect 7423 20825 7432 20859
rect 7380 20816 7432 20825
rect 9588 21088 9640 21140
rect 11336 21131 11388 21140
rect 11336 21097 11345 21131
rect 11345 21097 11379 21131
rect 11379 21097 11388 21131
rect 11336 21088 11388 21097
rect 12716 21088 12768 21140
rect 16212 21131 16264 21140
rect 16212 21097 16221 21131
rect 16221 21097 16255 21131
rect 16255 21097 16264 21131
rect 16212 21088 16264 21097
rect 18420 21131 18472 21140
rect 18420 21097 18429 21131
rect 18429 21097 18463 21131
rect 18463 21097 18472 21131
rect 18420 21088 18472 21097
rect 22284 21088 22336 21140
rect 23664 21088 23716 21140
rect 8944 20995 8996 21004
rect 8944 20961 8953 20995
rect 8953 20961 8987 20995
rect 8987 20961 8996 20995
rect 8944 20952 8996 20961
rect 14096 20995 14148 21004
rect 14096 20961 14105 20995
rect 14105 20961 14139 20995
rect 14139 20961 14148 20995
rect 14096 20952 14148 20961
rect 15384 20952 15436 21004
rect 15844 20952 15896 21004
rect 21272 21020 21324 21072
rect 8484 20884 8536 20936
rect 11888 20884 11940 20936
rect 12900 20884 12952 20936
rect 13820 20884 13872 20936
rect 16672 20927 16724 20936
rect 4804 20748 4856 20800
rect 7564 20791 7616 20800
rect 7564 20757 7589 20791
rect 7589 20757 7616 20791
rect 7564 20748 7616 20757
rect 9036 20748 9088 20800
rect 10416 20816 10468 20868
rect 14096 20816 14148 20868
rect 14740 20816 14792 20868
rect 16672 20893 16681 20927
rect 16681 20893 16715 20927
rect 16715 20893 16724 20927
rect 16672 20884 16724 20893
rect 16764 20927 16816 20936
rect 16764 20893 16773 20927
rect 16773 20893 16807 20927
rect 16807 20893 16816 20927
rect 17776 20927 17828 20936
rect 16764 20884 16816 20893
rect 16580 20816 16632 20868
rect 17776 20893 17785 20927
rect 17785 20893 17819 20927
rect 17819 20893 17828 20927
rect 17776 20884 17828 20893
rect 19432 20884 19484 20936
rect 25136 21088 25188 21140
rect 25320 21088 25372 21140
rect 24676 21020 24728 21072
rect 26976 21020 27028 21072
rect 27712 21020 27764 21072
rect 30288 21088 30340 21140
rect 31760 21088 31812 21140
rect 31944 21131 31996 21140
rect 31944 21097 31953 21131
rect 31953 21097 31987 21131
rect 31987 21097 31996 21131
rect 31944 21088 31996 21097
rect 34152 21088 34204 21140
rect 25136 20952 25188 21004
rect 24400 20927 24452 20936
rect 13820 20748 13872 20800
rect 18236 20816 18288 20868
rect 22652 20816 22704 20868
rect 23296 20859 23348 20868
rect 23296 20825 23305 20859
rect 23305 20825 23339 20859
rect 23339 20825 23348 20859
rect 23296 20816 23348 20825
rect 17224 20748 17276 20800
rect 18328 20748 18380 20800
rect 18696 20748 18748 20800
rect 19248 20748 19300 20800
rect 19432 20748 19484 20800
rect 24400 20893 24409 20927
rect 24409 20893 24443 20927
rect 24443 20893 24452 20927
rect 24400 20884 24452 20893
rect 24308 20816 24360 20868
rect 24584 20884 24636 20936
rect 26516 20884 26568 20936
rect 28172 20952 28224 21004
rect 29000 20884 29052 20936
rect 29828 20952 29880 21004
rect 30564 20927 30616 20936
rect 30564 20893 30573 20927
rect 30573 20893 30607 20927
rect 30607 20893 30616 20927
rect 30564 20884 30616 20893
rect 24676 20859 24728 20868
rect 24676 20825 24685 20859
rect 24685 20825 24719 20859
rect 24719 20825 24728 20859
rect 24676 20816 24728 20825
rect 25780 20816 25832 20868
rect 27068 20859 27120 20868
rect 27068 20825 27077 20859
rect 27077 20825 27111 20859
rect 27111 20825 27120 20859
rect 27068 20816 27120 20825
rect 24584 20748 24636 20800
rect 25688 20791 25740 20800
rect 25688 20757 25697 20791
rect 25697 20757 25731 20791
rect 25731 20757 25740 20791
rect 25688 20748 25740 20757
rect 26608 20748 26660 20800
rect 28080 20816 28132 20868
rect 30104 20816 30156 20868
rect 33508 20816 33560 20868
rect 33784 20859 33836 20868
rect 33784 20825 33793 20859
rect 33793 20825 33827 20859
rect 33827 20825 33836 20859
rect 33784 20816 33836 20825
rect 28448 20748 28500 20800
rect 28724 20748 28776 20800
rect 29828 20748 29880 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 5540 20587 5592 20596
rect 5540 20553 5565 20587
rect 5565 20553 5592 20587
rect 5724 20587 5776 20596
rect 5540 20544 5592 20553
rect 5724 20553 5733 20587
rect 5733 20553 5767 20587
rect 5767 20553 5776 20587
rect 5724 20544 5776 20553
rect 4620 20476 4672 20528
rect 5448 20476 5500 20528
rect 10416 20587 10468 20596
rect 5908 20476 5960 20528
rect 6460 20476 6512 20528
rect 10416 20553 10425 20587
rect 10425 20553 10459 20587
rect 10459 20553 10468 20587
rect 10416 20544 10468 20553
rect 12900 20544 12952 20596
rect 13912 20544 13964 20596
rect 14372 20544 14424 20596
rect 14740 20587 14792 20596
rect 14740 20553 14749 20587
rect 14749 20553 14783 20587
rect 14783 20553 14792 20587
rect 14740 20544 14792 20553
rect 15292 20544 15344 20596
rect 15660 20544 15712 20596
rect 7380 20519 7432 20528
rect 7380 20485 7389 20519
rect 7389 20485 7423 20519
rect 7423 20485 7432 20519
rect 7380 20476 7432 20485
rect 7564 20519 7616 20528
rect 7564 20485 7589 20519
rect 7589 20485 7616 20519
rect 7564 20476 7616 20485
rect 8944 20476 8996 20528
rect 16856 20519 16908 20528
rect 8668 20408 8720 20460
rect 9588 20408 9640 20460
rect 11520 20451 11572 20460
rect 11520 20417 11529 20451
rect 11529 20417 11563 20451
rect 11563 20417 11572 20451
rect 11520 20408 11572 20417
rect 13820 20408 13872 20460
rect 14648 20408 14700 20460
rect 14924 20451 14976 20460
rect 14924 20417 14933 20451
rect 14933 20417 14967 20451
rect 14967 20417 14976 20451
rect 14924 20408 14976 20417
rect 15108 20408 15160 20460
rect 2872 20247 2924 20256
rect 2872 20213 2881 20247
rect 2881 20213 2915 20247
rect 2915 20213 2924 20247
rect 2872 20204 2924 20213
rect 3792 20204 3844 20256
rect 6552 20247 6604 20256
rect 6552 20213 6561 20247
rect 6561 20213 6595 20247
rect 6595 20213 6604 20247
rect 6552 20204 6604 20213
rect 8392 20204 8444 20256
rect 15568 20408 15620 20460
rect 16856 20485 16865 20519
rect 16865 20485 16899 20519
rect 16899 20485 16908 20519
rect 16856 20476 16908 20485
rect 17776 20544 17828 20596
rect 20076 20544 20128 20596
rect 25412 20544 25464 20596
rect 16488 20408 16540 20460
rect 16764 20408 16816 20460
rect 17960 20451 18012 20460
rect 17960 20417 17969 20451
rect 17969 20417 18003 20451
rect 18003 20417 18012 20451
rect 18144 20451 18196 20460
rect 17960 20408 18012 20417
rect 18144 20417 18153 20451
rect 18153 20417 18187 20451
rect 18187 20417 18196 20451
rect 18144 20408 18196 20417
rect 18236 20451 18288 20460
rect 18236 20417 18245 20451
rect 18245 20417 18279 20451
rect 18279 20417 18288 20451
rect 18788 20476 18840 20528
rect 18236 20408 18288 20417
rect 20076 20451 20128 20460
rect 20076 20417 20085 20451
rect 20085 20417 20119 20451
rect 20119 20417 20128 20451
rect 20076 20408 20128 20417
rect 18328 20340 18380 20392
rect 16672 20272 16724 20324
rect 16028 20204 16080 20256
rect 16580 20204 16632 20256
rect 17040 20247 17092 20256
rect 17040 20213 17049 20247
rect 17049 20213 17083 20247
rect 17083 20213 17092 20247
rect 17040 20204 17092 20213
rect 18420 20204 18472 20256
rect 20076 20272 20128 20324
rect 20260 20451 20312 20460
rect 20260 20417 20269 20451
rect 20269 20417 20303 20451
rect 20303 20417 20312 20451
rect 20444 20451 20496 20460
rect 20260 20408 20312 20417
rect 20444 20417 20453 20451
rect 20453 20417 20487 20451
rect 20487 20417 20496 20451
rect 20444 20408 20496 20417
rect 20904 20476 20956 20528
rect 22008 20408 22060 20460
rect 23572 20476 23624 20528
rect 24492 20451 24544 20460
rect 24492 20417 24501 20451
rect 24501 20417 24535 20451
rect 24535 20417 24544 20451
rect 24492 20408 24544 20417
rect 25136 20451 25188 20460
rect 24124 20340 24176 20392
rect 24308 20340 24360 20392
rect 25136 20417 25145 20451
rect 25145 20417 25179 20451
rect 25179 20417 25188 20451
rect 25136 20408 25188 20417
rect 25228 20451 25280 20460
rect 25228 20417 25238 20451
rect 25238 20417 25272 20451
rect 25272 20417 25280 20451
rect 25412 20451 25464 20460
rect 25228 20408 25280 20417
rect 25412 20417 25421 20451
rect 25421 20417 25455 20451
rect 25455 20417 25464 20451
rect 25412 20408 25464 20417
rect 26884 20544 26936 20596
rect 27252 20476 27304 20528
rect 27804 20544 27856 20596
rect 28724 20544 28776 20596
rect 28816 20544 28868 20596
rect 29000 20544 29052 20596
rect 29920 20544 29972 20596
rect 30196 20544 30248 20596
rect 28356 20476 28408 20528
rect 27804 20451 27856 20460
rect 24860 20340 24912 20392
rect 27804 20417 27813 20451
rect 27813 20417 27847 20451
rect 27847 20417 27856 20451
rect 27804 20408 27856 20417
rect 28080 20408 28132 20460
rect 29828 20519 29880 20528
rect 29828 20485 29862 20519
rect 29862 20485 29880 20519
rect 29828 20476 29880 20485
rect 26700 20340 26752 20392
rect 28908 20451 28960 20460
rect 28908 20417 28917 20451
rect 28917 20417 28951 20451
rect 28951 20417 28960 20451
rect 28908 20408 28960 20417
rect 30748 20408 30800 20460
rect 31760 20408 31812 20460
rect 33876 20408 33928 20460
rect 34520 20408 34572 20460
rect 29368 20340 29420 20392
rect 21732 20272 21784 20324
rect 21088 20204 21140 20256
rect 23480 20204 23532 20256
rect 23756 20204 23808 20256
rect 24676 20204 24728 20256
rect 26516 20204 26568 20256
rect 26976 20204 27028 20256
rect 28724 20272 28776 20324
rect 33692 20340 33744 20392
rect 34796 20340 34848 20392
rect 31300 20272 31352 20324
rect 32864 20272 32916 20324
rect 29000 20204 29052 20256
rect 29368 20204 29420 20256
rect 30932 20247 30984 20256
rect 30932 20213 30941 20247
rect 30941 20213 30975 20247
rect 30975 20213 30984 20247
rect 30932 20204 30984 20213
rect 32312 20247 32364 20256
rect 32312 20213 32321 20247
rect 32321 20213 32355 20247
rect 32355 20213 32364 20247
rect 32312 20204 32364 20213
rect 33140 20204 33192 20256
rect 34336 20204 34388 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 6552 20000 6604 20052
rect 2872 19864 2924 19916
rect 8668 20000 8720 20052
rect 8484 19932 8536 19984
rect 17316 20000 17368 20052
rect 14556 19932 14608 19984
rect 15568 19932 15620 19984
rect 18328 19932 18380 19984
rect 8944 19907 8996 19916
rect 3792 19839 3844 19848
rect 3792 19805 3801 19839
rect 3801 19805 3835 19839
rect 3835 19805 3844 19839
rect 3792 19796 3844 19805
rect 8944 19873 8953 19907
rect 8953 19873 8987 19907
rect 8987 19873 8996 19907
rect 8944 19864 8996 19873
rect 6920 19839 6972 19848
rect 6920 19805 6929 19839
rect 6929 19805 6963 19839
rect 6963 19805 6972 19839
rect 6920 19796 6972 19805
rect 8392 19839 8444 19848
rect 8392 19805 8401 19839
rect 8401 19805 8435 19839
rect 8435 19805 8444 19839
rect 8392 19796 8444 19805
rect 9036 19796 9088 19848
rect 10876 19796 10928 19848
rect 15200 19796 15252 19848
rect 7380 19771 7432 19780
rect 7380 19737 7389 19771
rect 7389 19737 7423 19771
rect 7423 19737 7432 19771
rect 7380 19728 7432 19737
rect 7564 19771 7616 19780
rect 7564 19737 7589 19771
rect 7589 19737 7616 19771
rect 7564 19728 7616 19737
rect 11060 19728 11112 19780
rect 11704 19728 11756 19780
rect 14004 19728 14056 19780
rect 14280 19771 14332 19780
rect 14280 19737 14289 19771
rect 14289 19737 14323 19771
rect 14323 19737 14332 19771
rect 14280 19728 14332 19737
rect 16304 19796 16356 19848
rect 18236 19839 18288 19848
rect 18236 19805 18245 19839
rect 18245 19805 18279 19839
rect 18279 19805 18288 19839
rect 18236 19796 18288 19805
rect 20628 20000 20680 20052
rect 20812 20000 20864 20052
rect 23388 20000 23440 20052
rect 21732 19907 21784 19916
rect 18420 19839 18472 19848
rect 18420 19805 18429 19839
rect 18429 19805 18463 19839
rect 18463 19805 18472 19839
rect 18420 19796 18472 19805
rect 18696 19796 18748 19848
rect 21732 19873 21741 19907
rect 21741 19873 21775 19907
rect 21775 19873 21784 19907
rect 21732 19864 21784 19873
rect 22008 19907 22060 19916
rect 22008 19873 22017 19907
rect 22017 19873 22051 19907
rect 22051 19873 22060 19907
rect 22008 19864 22060 19873
rect 23204 19864 23256 19916
rect 20444 19796 20496 19848
rect 22652 19796 22704 19848
rect 23572 19864 23624 19916
rect 23480 19839 23532 19848
rect 23480 19805 23489 19839
rect 23489 19805 23523 19839
rect 23523 19805 23532 19839
rect 25228 20000 25280 20052
rect 30564 20000 30616 20052
rect 33692 20043 33744 20052
rect 25136 19932 25188 19984
rect 24676 19864 24728 19916
rect 23480 19796 23532 19805
rect 24492 19839 24544 19848
rect 24492 19805 24502 19839
rect 24502 19805 24536 19839
rect 24536 19805 24544 19839
rect 24492 19796 24544 19805
rect 6460 19660 6512 19712
rect 12348 19703 12400 19712
rect 12348 19669 12357 19703
rect 12357 19669 12391 19703
rect 12391 19669 12400 19703
rect 12348 19660 12400 19669
rect 13820 19660 13872 19712
rect 16396 19728 16448 19780
rect 16764 19728 16816 19780
rect 20168 19771 20220 19780
rect 20168 19737 20202 19771
rect 20202 19737 20220 19771
rect 20168 19728 20220 19737
rect 23756 19728 23808 19780
rect 24860 19839 24912 19848
rect 24860 19805 24874 19839
rect 24874 19805 24908 19839
rect 24908 19805 24912 19839
rect 24860 19796 24912 19805
rect 25136 19796 25188 19848
rect 26700 19839 26752 19848
rect 15200 19703 15252 19712
rect 15200 19669 15209 19703
rect 15209 19669 15243 19703
rect 15243 19669 15252 19703
rect 15200 19660 15252 19669
rect 16580 19660 16632 19712
rect 18420 19660 18472 19712
rect 22376 19660 22428 19712
rect 23020 19703 23072 19712
rect 23020 19669 23029 19703
rect 23029 19669 23063 19703
rect 23063 19669 23072 19703
rect 23020 19660 23072 19669
rect 25412 19728 25464 19780
rect 24952 19660 25004 19712
rect 26700 19805 26709 19839
rect 26709 19805 26743 19839
rect 26743 19805 26752 19839
rect 26700 19796 26752 19805
rect 26884 19796 26936 19848
rect 27436 19796 27488 19848
rect 27712 19932 27764 19984
rect 28172 19932 28224 19984
rect 29000 19932 29052 19984
rect 31300 19932 31352 19984
rect 28448 19864 28500 19916
rect 33692 20009 33701 20043
rect 33701 20009 33735 20043
rect 33735 20009 33744 20043
rect 33692 20000 33744 20009
rect 27896 19839 27948 19848
rect 27896 19805 27905 19839
rect 27905 19805 27939 19839
rect 27939 19805 27948 19839
rect 27896 19796 27948 19805
rect 28172 19796 28224 19848
rect 33784 19864 33836 19916
rect 32956 19796 33008 19848
rect 28356 19728 28408 19780
rect 32220 19728 32272 19780
rect 26700 19660 26752 19712
rect 27160 19660 27212 19712
rect 27436 19703 27488 19712
rect 27436 19669 27445 19703
rect 27445 19669 27479 19703
rect 27479 19669 27488 19703
rect 27436 19660 27488 19669
rect 37280 19660 37332 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 5080 19456 5132 19508
rect 5356 19388 5408 19440
rect 5540 19388 5592 19440
rect 9496 19456 9548 19508
rect 10876 19456 10928 19508
rect 5632 19320 5684 19372
rect 5816 19363 5868 19372
rect 5816 19329 5825 19363
rect 5825 19329 5859 19363
rect 5859 19329 5868 19363
rect 5816 19320 5868 19329
rect 8944 19388 8996 19440
rect 9220 19388 9272 19440
rect 8668 19320 8720 19372
rect 10784 19363 10836 19372
rect 10784 19329 10793 19363
rect 10793 19329 10827 19363
rect 10827 19329 10836 19363
rect 10784 19320 10836 19329
rect 14280 19456 14332 19508
rect 16764 19456 16816 19508
rect 17132 19456 17184 19508
rect 20444 19499 20496 19508
rect 15200 19388 15252 19440
rect 15936 19363 15988 19372
rect 15936 19329 15945 19363
rect 15945 19329 15979 19363
rect 15979 19329 15988 19363
rect 15936 19320 15988 19329
rect 16028 19320 16080 19372
rect 11704 19252 11756 19304
rect 17960 19388 18012 19440
rect 18236 19388 18288 19440
rect 18972 19388 19024 19440
rect 17316 19363 17368 19372
rect 17316 19329 17325 19363
rect 17325 19329 17359 19363
rect 17359 19329 17368 19363
rect 17316 19320 17368 19329
rect 17868 19320 17920 19372
rect 20444 19465 20453 19499
rect 20453 19465 20487 19499
rect 20487 19465 20496 19499
rect 20444 19456 20496 19465
rect 24032 19456 24084 19508
rect 24768 19456 24820 19508
rect 23020 19388 23072 19440
rect 20444 19320 20496 19372
rect 19432 19252 19484 19304
rect 16672 19227 16724 19236
rect 16672 19193 16681 19227
rect 16681 19193 16715 19227
rect 16715 19193 16724 19227
rect 16672 19184 16724 19193
rect 23756 19320 23808 19372
rect 24860 19388 24912 19440
rect 25044 19388 25096 19440
rect 26700 19388 26752 19440
rect 27804 19456 27856 19508
rect 30196 19499 30248 19508
rect 30196 19465 30205 19499
rect 30205 19465 30239 19499
rect 30239 19465 30248 19499
rect 30196 19456 30248 19465
rect 32220 19499 32272 19508
rect 32220 19465 32229 19499
rect 32229 19465 32263 19499
rect 32263 19465 32272 19499
rect 32220 19456 32272 19465
rect 34704 19456 34756 19508
rect 34796 19456 34848 19508
rect 27436 19388 27488 19440
rect 24400 19363 24452 19372
rect 24400 19329 24434 19363
rect 24434 19329 24452 19363
rect 24400 19320 24452 19329
rect 27068 19320 27120 19372
rect 28816 19363 28868 19372
rect 28816 19329 28825 19363
rect 28825 19329 28859 19363
rect 28859 19329 28868 19363
rect 28816 19320 28868 19329
rect 30840 19320 30892 19372
rect 32404 19363 32456 19372
rect 32404 19329 32413 19363
rect 32413 19329 32447 19363
rect 32447 19329 32456 19363
rect 32404 19320 32456 19329
rect 33140 19363 33192 19372
rect 33140 19329 33149 19363
rect 33149 19329 33183 19363
rect 33183 19329 33192 19363
rect 33140 19320 33192 19329
rect 33600 19320 33652 19372
rect 34428 19388 34480 19440
rect 34336 19320 34388 19372
rect 37648 19320 37700 19372
rect 32956 19295 33008 19304
rect 32956 19261 32965 19295
rect 32965 19261 32999 19295
rect 32999 19261 33008 19295
rect 32956 19252 33008 19261
rect 37280 19295 37332 19304
rect 37280 19261 37289 19295
rect 37289 19261 37323 19295
rect 37323 19261 37332 19295
rect 37280 19252 37332 19261
rect 4804 19159 4856 19168
rect 4804 19125 4813 19159
rect 4813 19125 4847 19159
rect 4847 19125 4856 19159
rect 4804 19116 4856 19125
rect 7748 19159 7800 19168
rect 7748 19125 7757 19159
rect 7757 19125 7791 19159
rect 7791 19125 7800 19159
rect 7748 19116 7800 19125
rect 11152 19116 11204 19168
rect 15200 19116 15252 19168
rect 24308 19116 24360 19168
rect 30748 19159 30800 19168
rect 30748 19125 30757 19159
rect 30757 19125 30791 19159
rect 30791 19125 30800 19159
rect 30748 19116 30800 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 3792 18912 3844 18964
rect 5540 18912 5592 18964
rect 7748 18912 7800 18964
rect 8668 18912 8720 18964
rect 11060 18912 11112 18964
rect 5816 18844 5868 18896
rect 8392 18776 8444 18828
rect 9220 18776 9272 18828
rect 8300 18751 8352 18760
rect 8300 18717 8309 18751
rect 8309 18717 8343 18751
rect 8343 18717 8352 18751
rect 8300 18708 8352 18717
rect 10508 18708 10560 18760
rect 6460 18683 6512 18692
rect 6460 18649 6469 18683
rect 6469 18649 6503 18683
rect 6503 18649 6512 18683
rect 6460 18640 6512 18649
rect 5356 18572 5408 18624
rect 11060 18708 11112 18760
rect 12624 18776 12676 18828
rect 12072 18751 12124 18760
rect 12072 18717 12081 18751
rect 12081 18717 12115 18751
rect 12115 18717 12124 18751
rect 12072 18708 12124 18717
rect 13176 18751 13228 18760
rect 13176 18717 13185 18751
rect 13185 18717 13219 18751
rect 13219 18717 13228 18751
rect 13176 18708 13228 18717
rect 15568 18844 15620 18896
rect 13820 18776 13872 18828
rect 14004 18776 14056 18828
rect 17592 18912 17644 18964
rect 15752 18844 15804 18896
rect 15752 18751 15804 18760
rect 15752 18717 15761 18751
rect 15761 18717 15795 18751
rect 15795 18717 15804 18751
rect 15752 18708 15804 18717
rect 19248 18844 19300 18896
rect 20904 18912 20956 18964
rect 24400 18955 24452 18964
rect 24400 18921 24409 18955
rect 24409 18921 24443 18955
rect 24443 18921 24452 18955
rect 24400 18912 24452 18921
rect 27068 18912 27120 18964
rect 27896 18912 27948 18964
rect 34520 18912 34572 18964
rect 16580 18776 16632 18828
rect 16212 18708 16264 18760
rect 16856 18751 16908 18760
rect 11980 18640 12032 18692
rect 14004 18640 14056 18692
rect 15016 18640 15068 18692
rect 16856 18717 16865 18751
rect 16865 18717 16899 18751
rect 16899 18717 16908 18751
rect 16856 18708 16908 18717
rect 10968 18572 11020 18624
rect 12256 18572 12308 18624
rect 12900 18615 12952 18624
rect 12900 18581 12909 18615
rect 12909 18581 12943 18615
rect 12943 18581 12952 18615
rect 12900 18572 12952 18581
rect 16304 18572 16356 18624
rect 16580 18615 16632 18624
rect 16580 18581 16589 18615
rect 16589 18581 16623 18615
rect 16623 18581 16632 18615
rect 16580 18572 16632 18581
rect 17040 18751 17092 18760
rect 17040 18717 17049 18751
rect 17049 18717 17083 18751
rect 17083 18717 17092 18751
rect 17040 18708 17092 18717
rect 18328 18751 18380 18760
rect 18328 18717 18337 18751
rect 18337 18717 18371 18751
rect 18371 18717 18380 18751
rect 18328 18708 18380 18717
rect 19340 18776 19392 18828
rect 21640 18844 21692 18896
rect 22100 18844 22152 18896
rect 23112 18844 23164 18896
rect 18604 18708 18656 18760
rect 18696 18751 18748 18760
rect 18696 18717 18705 18751
rect 18705 18717 18739 18751
rect 18739 18717 18748 18751
rect 18696 18708 18748 18717
rect 21447 18748 21499 18760
rect 21447 18714 21480 18748
rect 21480 18714 21499 18748
rect 19984 18640 20036 18692
rect 21447 18708 21499 18714
rect 20352 18640 20404 18692
rect 22008 18708 22060 18760
rect 17224 18572 17276 18624
rect 19064 18572 19116 18624
rect 21180 18572 21232 18624
rect 23572 18776 23624 18828
rect 27344 18844 27396 18896
rect 22376 18751 22428 18760
rect 22376 18717 22385 18751
rect 22385 18717 22419 18751
rect 22419 18717 22428 18751
rect 22376 18708 22428 18717
rect 23296 18708 23348 18760
rect 23204 18640 23256 18692
rect 23388 18572 23440 18624
rect 24492 18640 24544 18692
rect 25228 18708 25280 18760
rect 26608 18708 26660 18760
rect 26976 18751 27028 18760
rect 26976 18717 26985 18751
rect 26985 18717 27019 18751
rect 27019 18717 27028 18751
rect 28172 18776 28224 18828
rect 32956 18776 33008 18828
rect 34704 18819 34756 18828
rect 34704 18785 34713 18819
rect 34713 18785 34747 18819
rect 34747 18785 34756 18819
rect 34704 18776 34756 18785
rect 26976 18708 27028 18717
rect 27252 18708 27304 18760
rect 28080 18708 28132 18760
rect 30656 18751 30708 18760
rect 30656 18717 30665 18751
rect 30665 18717 30699 18751
rect 30699 18717 30708 18751
rect 30656 18708 30708 18717
rect 30748 18708 30800 18760
rect 32772 18751 32824 18760
rect 32772 18717 32781 18751
rect 32781 18717 32815 18751
rect 32815 18717 32824 18751
rect 32772 18708 32824 18717
rect 33140 18708 33192 18760
rect 34980 18751 35032 18760
rect 34980 18717 34989 18751
rect 34989 18717 35023 18751
rect 35023 18717 35032 18751
rect 34980 18708 35032 18717
rect 33692 18683 33744 18692
rect 33692 18649 33701 18683
rect 33701 18649 33735 18683
rect 33735 18649 33744 18683
rect 33692 18640 33744 18649
rect 25228 18572 25280 18624
rect 30932 18572 30984 18624
rect 33048 18572 33100 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 6920 18368 6972 18420
rect 10784 18368 10836 18420
rect 11980 18368 12032 18420
rect 14648 18368 14700 18420
rect 14924 18368 14976 18420
rect 12348 18300 12400 18352
rect 17868 18368 17920 18420
rect 8852 18232 8904 18284
rect 8944 18232 8996 18284
rect 11612 18232 11664 18284
rect 11704 18275 11756 18284
rect 11704 18241 11713 18275
rect 11713 18241 11747 18275
rect 11747 18241 11756 18275
rect 11704 18232 11756 18241
rect 13084 18232 13136 18284
rect 14556 18232 14608 18284
rect 15200 18300 15252 18352
rect 16396 18300 16448 18352
rect 15016 18275 15068 18284
rect 15016 18241 15025 18275
rect 15025 18241 15059 18275
rect 15059 18241 15068 18275
rect 15016 18232 15068 18241
rect 16028 18232 16080 18284
rect 17224 18232 17276 18284
rect 17592 18275 17644 18284
rect 17592 18241 17601 18275
rect 17601 18241 17635 18275
rect 17635 18241 17644 18275
rect 17592 18232 17644 18241
rect 19340 18300 19392 18352
rect 10968 18096 11020 18148
rect 14924 18096 14976 18148
rect 15108 18096 15160 18148
rect 18604 18275 18656 18284
rect 18604 18241 18613 18275
rect 18613 18241 18647 18275
rect 18647 18241 18656 18275
rect 18604 18232 18656 18241
rect 20168 18368 20220 18420
rect 23112 18343 23164 18352
rect 19892 18232 19944 18284
rect 19616 18164 19668 18216
rect 14372 18071 14424 18080
rect 14372 18037 14381 18071
rect 14381 18037 14415 18071
rect 14415 18037 14424 18071
rect 14372 18028 14424 18037
rect 14740 18028 14792 18080
rect 15752 18028 15804 18080
rect 18604 18096 18656 18148
rect 19708 18096 19760 18148
rect 20352 18275 20404 18284
rect 20352 18241 20361 18275
rect 20361 18241 20395 18275
rect 20395 18241 20404 18275
rect 20352 18232 20404 18241
rect 20812 18232 20864 18284
rect 23112 18309 23121 18343
rect 23121 18309 23155 18343
rect 23155 18309 23164 18343
rect 23112 18300 23164 18309
rect 24308 18343 24360 18352
rect 24308 18309 24317 18343
rect 24317 18309 24351 18343
rect 24351 18309 24360 18343
rect 24308 18300 24360 18309
rect 32404 18368 32456 18420
rect 25044 18300 25096 18352
rect 25596 18300 25648 18352
rect 32312 18343 32364 18352
rect 32312 18309 32321 18343
rect 32321 18309 32355 18343
rect 32355 18309 32364 18343
rect 32312 18300 32364 18309
rect 21640 18232 21692 18284
rect 21916 18232 21968 18284
rect 22560 18232 22612 18284
rect 23388 18232 23440 18284
rect 24124 18275 24176 18284
rect 24124 18241 24133 18275
rect 24133 18241 24167 18275
rect 24167 18241 24176 18275
rect 24124 18232 24176 18241
rect 27252 18232 27304 18284
rect 30472 18232 30524 18284
rect 30932 18275 30984 18284
rect 30932 18241 30941 18275
rect 30941 18241 30975 18275
rect 30975 18241 30984 18275
rect 30932 18232 30984 18241
rect 32128 18275 32180 18284
rect 32128 18241 32137 18275
rect 32137 18241 32171 18275
rect 32171 18241 32180 18275
rect 32128 18232 32180 18241
rect 33048 18275 33100 18284
rect 33048 18241 33057 18275
rect 33057 18241 33091 18275
rect 33091 18241 33100 18275
rect 33048 18232 33100 18241
rect 21456 18164 21508 18216
rect 20904 18096 20956 18148
rect 21272 18096 21324 18148
rect 24492 18139 24544 18148
rect 24492 18105 24501 18139
rect 24501 18105 24535 18139
rect 24535 18105 24544 18139
rect 24492 18096 24544 18105
rect 24676 18096 24728 18148
rect 32956 18164 33008 18216
rect 33508 18164 33560 18216
rect 34520 18164 34572 18216
rect 37832 18164 37884 18216
rect 21732 18028 21784 18080
rect 22008 18028 22060 18080
rect 23296 18028 23348 18080
rect 25136 18028 25188 18080
rect 30564 18028 30616 18080
rect 30748 18028 30800 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 8852 17824 8904 17876
rect 5908 17756 5960 17808
rect 9404 17756 9456 17808
rect 11520 17824 11572 17876
rect 11612 17824 11664 17876
rect 13176 17824 13228 17876
rect 14556 17824 14608 17876
rect 16856 17824 16908 17876
rect 19616 17867 19668 17876
rect 19616 17833 19625 17867
rect 19625 17833 19659 17867
rect 19659 17833 19668 17867
rect 19616 17824 19668 17833
rect 11152 17756 11204 17808
rect 5816 17620 5868 17672
rect 7104 17663 7156 17672
rect 7104 17629 7113 17663
rect 7113 17629 7147 17663
rect 7147 17629 7156 17663
rect 7104 17620 7156 17629
rect 10968 17663 11020 17672
rect 10968 17629 10977 17663
rect 10977 17629 11011 17663
rect 11011 17629 11020 17663
rect 10968 17620 11020 17629
rect 11152 17663 11204 17672
rect 11152 17629 11161 17663
rect 11161 17629 11195 17663
rect 11195 17629 11204 17663
rect 11336 17663 11388 17672
rect 11152 17620 11204 17629
rect 11336 17629 11345 17663
rect 11345 17629 11379 17663
rect 11379 17629 11388 17663
rect 11336 17620 11388 17629
rect 11980 17620 12032 17672
rect 15292 17756 15344 17808
rect 12808 17688 12860 17740
rect 13452 17688 13504 17740
rect 20720 17824 20772 17876
rect 22560 17867 22612 17876
rect 22560 17833 22569 17867
rect 22569 17833 22603 17867
rect 22603 17833 22612 17867
rect 22560 17824 22612 17833
rect 23296 17824 23348 17876
rect 30840 17867 30892 17876
rect 20444 17756 20496 17808
rect 24860 17731 24912 17740
rect 24860 17697 24869 17731
rect 24869 17697 24903 17731
rect 24903 17697 24912 17731
rect 24860 17688 24912 17697
rect 28172 17688 28224 17740
rect 28632 17731 28684 17740
rect 28632 17697 28641 17731
rect 28641 17697 28675 17731
rect 28675 17697 28684 17731
rect 28632 17688 28684 17697
rect 30840 17833 30849 17867
rect 30849 17833 30883 17867
rect 30883 17833 30892 17867
rect 30840 17824 30892 17833
rect 34520 17824 34572 17876
rect 32128 17688 32180 17740
rect 32312 17688 32364 17740
rect 9404 17595 9456 17604
rect 9404 17561 9413 17595
rect 9413 17561 9447 17595
rect 9447 17561 9456 17595
rect 9404 17552 9456 17561
rect 12624 17620 12676 17672
rect 13820 17620 13872 17672
rect 15476 17620 15528 17672
rect 17592 17620 17644 17672
rect 19432 17663 19484 17672
rect 19432 17629 19441 17663
rect 19441 17629 19475 17663
rect 19475 17629 19484 17663
rect 19432 17620 19484 17629
rect 20076 17620 20128 17672
rect 15016 17595 15068 17604
rect 15016 17561 15025 17595
rect 15025 17561 15059 17595
rect 15059 17561 15068 17595
rect 15016 17552 15068 17561
rect 16028 17552 16080 17604
rect 17224 17595 17276 17604
rect 17224 17561 17233 17595
rect 17233 17561 17267 17595
rect 17267 17561 17276 17595
rect 17224 17552 17276 17561
rect 19340 17552 19392 17604
rect 6184 17484 6236 17536
rect 9956 17484 10008 17536
rect 12072 17484 12124 17536
rect 13084 17484 13136 17536
rect 16212 17484 16264 17536
rect 17132 17484 17184 17536
rect 20352 17484 20404 17536
rect 20720 17663 20772 17672
rect 20720 17629 20729 17663
rect 20729 17629 20763 17663
rect 20763 17629 20772 17663
rect 20720 17620 20772 17629
rect 21732 17620 21784 17672
rect 23204 17663 23256 17672
rect 23204 17629 23213 17663
rect 23213 17629 23247 17663
rect 23247 17629 23256 17663
rect 23204 17620 23256 17629
rect 28356 17663 28408 17672
rect 28356 17629 28365 17663
rect 28365 17629 28399 17663
rect 28399 17629 28408 17663
rect 28356 17620 28408 17629
rect 21272 17552 21324 17604
rect 22468 17552 22520 17604
rect 26976 17552 27028 17604
rect 30564 17552 30616 17604
rect 32956 17620 33008 17672
rect 34428 17620 34480 17672
rect 33692 17552 33744 17604
rect 21640 17484 21692 17536
rect 22560 17484 22612 17536
rect 26148 17484 26200 17536
rect 28908 17484 28960 17536
rect 29920 17484 29972 17536
rect 30472 17484 30524 17536
rect 33140 17484 33192 17536
rect 36084 17527 36136 17536
rect 36084 17493 36093 17527
rect 36093 17493 36127 17527
rect 36127 17493 36136 17527
rect 36084 17484 36136 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 4068 17280 4120 17332
rect 12532 17323 12584 17332
rect 12532 17289 12541 17323
rect 12541 17289 12575 17323
rect 12575 17289 12584 17323
rect 12532 17280 12584 17289
rect 12992 17280 13044 17332
rect 13452 17323 13504 17332
rect 13452 17289 13461 17323
rect 13461 17289 13495 17323
rect 13495 17289 13504 17323
rect 13452 17280 13504 17289
rect 15016 17280 15068 17332
rect 18696 17280 18748 17332
rect 6092 17212 6144 17264
rect 5448 17144 5500 17196
rect 2688 17119 2740 17128
rect 2688 17085 2697 17119
rect 2697 17085 2731 17119
rect 2731 17085 2740 17119
rect 2688 17076 2740 17085
rect 3700 17076 3752 17128
rect 7012 17144 7064 17196
rect 7380 17187 7432 17196
rect 7380 17153 7389 17187
rect 7389 17153 7423 17187
rect 7423 17153 7432 17187
rect 7380 17144 7432 17153
rect 13084 17212 13136 17264
rect 9312 17144 9364 17196
rect 4620 17008 4672 17060
rect 8116 17076 8168 17128
rect 8852 17076 8904 17128
rect 13820 17144 13872 17196
rect 15752 17212 15804 17264
rect 16028 17212 16080 17264
rect 14280 17144 14332 17196
rect 15016 17144 15068 17196
rect 15384 17187 15436 17196
rect 14556 17076 14608 17128
rect 15384 17153 15393 17187
rect 15393 17153 15427 17187
rect 15427 17153 15436 17187
rect 15384 17144 15436 17153
rect 15476 17187 15528 17196
rect 15476 17153 15485 17187
rect 15485 17153 15519 17187
rect 15519 17153 15528 17187
rect 15936 17187 15988 17196
rect 15476 17144 15528 17153
rect 15936 17153 15945 17187
rect 15945 17153 15979 17187
rect 15979 17153 15988 17187
rect 15936 17144 15988 17153
rect 17868 17144 17920 17196
rect 19524 17144 19576 17196
rect 20076 17280 20128 17332
rect 20812 17280 20864 17332
rect 20536 17212 20588 17264
rect 15568 17076 15620 17128
rect 17224 17076 17276 17128
rect 12624 17008 12676 17060
rect 15752 17008 15804 17060
rect 18604 17076 18656 17128
rect 19432 17119 19484 17128
rect 19432 17085 19441 17119
rect 19441 17085 19475 17119
rect 19475 17085 19484 17119
rect 19432 17076 19484 17085
rect 20168 17144 20220 17196
rect 22468 17280 22520 17332
rect 26976 17323 27028 17332
rect 26976 17289 26985 17323
rect 26985 17289 27019 17323
rect 27019 17289 27028 17323
rect 26976 17280 27028 17289
rect 28356 17280 28408 17332
rect 31852 17280 31904 17332
rect 20720 17076 20772 17128
rect 5540 16940 5592 16992
rect 8208 16940 8260 16992
rect 14924 16983 14976 16992
rect 14924 16949 14933 16983
rect 14933 16949 14967 16983
rect 14967 16949 14976 16983
rect 14924 16940 14976 16949
rect 16028 16983 16080 16992
rect 16028 16949 16037 16983
rect 16037 16949 16071 16983
rect 16071 16949 16080 16983
rect 16028 16940 16080 16949
rect 17040 16940 17092 16992
rect 19248 17008 19300 17060
rect 20168 17008 20220 17060
rect 21456 17144 21508 17196
rect 23296 17187 23348 17196
rect 23296 17153 23305 17187
rect 23305 17153 23339 17187
rect 23339 17153 23348 17187
rect 23296 17144 23348 17153
rect 24676 17144 24728 17196
rect 25596 17144 25648 17196
rect 26148 17187 26200 17196
rect 21640 17076 21692 17128
rect 22376 17076 22428 17128
rect 26148 17153 26157 17187
rect 26157 17153 26191 17187
rect 26191 17153 26200 17187
rect 26148 17144 26200 17153
rect 26332 17076 26384 17128
rect 27252 17076 27304 17128
rect 28816 17212 28868 17264
rect 28632 17144 28684 17196
rect 30656 17212 30708 17264
rect 33416 17212 33468 17264
rect 29828 17144 29880 17196
rect 31300 17144 31352 17196
rect 34152 17212 34204 17264
rect 31944 17076 31996 17128
rect 34428 17076 34480 17128
rect 25044 17008 25096 17060
rect 26148 17008 26200 17060
rect 33968 17008 34020 17060
rect 20076 16940 20128 16992
rect 20536 16983 20588 16992
rect 20536 16949 20545 16983
rect 20545 16949 20579 16983
rect 20579 16949 20588 16983
rect 20536 16940 20588 16949
rect 25596 16940 25648 16992
rect 30840 16940 30892 16992
rect 32496 16983 32548 16992
rect 32496 16949 32505 16983
rect 32505 16949 32539 16983
rect 32539 16949 32548 16983
rect 32496 16940 32548 16949
rect 33784 16940 33836 16992
rect 34520 16940 34572 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 7380 16779 7432 16788
rect 7380 16745 7389 16779
rect 7389 16745 7423 16779
rect 7423 16745 7432 16779
rect 7380 16736 7432 16745
rect 9036 16736 9088 16788
rect 9312 16779 9364 16788
rect 9312 16745 9321 16779
rect 9321 16745 9355 16779
rect 9355 16745 9364 16779
rect 9312 16736 9364 16745
rect 2872 16600 2924 16652
rect 3792 16643 3844 16652
rect 3792 16609 3801 16643
rect 3801 16609 3835 16643
rect 3835 16609 3844 16643
rect 3792 16600 3844 16609
rect 1860 16575 1912 16584
rect 1860 16541 1869 16575
rect 1869 16541 1903 16575
rect 1903 16541 1912 16575
rect 1860 16532 1912 16541
rect 2688 16532 2740 16584
rect 4068 16575 4120 16584
rect 4068 16541 4102 16575
rect 4102 16541 4120 16575
rect 4068 16532 4120 16541
rect 8852 16668 8904 16720
rect 10692 16668 10744 16720
rect 13728 16736 13780 16788
rect 15016 16736 15068 16788
rect 5724 16464 5776 16516
rect 6000 16464 6052 16516
rect 7012 16507 7064 16516
rect 5080 16396 5132 16448
rect 5632 16396 5684 16448
rect 7012 16473 7021 16507
rect 7021 16473 7055 16507
rect 7055 16473 7064 16507
rect 7012 16464 7064 16473
rect 7196 16396 7248 16448
rect 10968 16532 11020 16584
rect 11336 16600 11388 16652
rect 11244 16575 11296 16584
rect 11244 16541 11258 16575
rect 11258 16541 11292 16575
rect 11292 16541 11296 16575
rect 11244 16532 11296 16541
rect 8944 16507 8996 16516
rect 8944 16473 8953 16507
rect 8953 16473 8987 16507
rect 8987 16473 8996 16507
rect 8944 16464 8996 16473
rect 9128 16507 9180 16516
rect 9128 16473 9137 16507
rect 9137 16473 9171 16507
rect 9171 16473 9180 16507
rect 9128 16464 9180 16473
rect 14740 16668 14792 16720
rect 13084 16532 13136 16584
rect 13268 16538 13274 16562
rect 13274 16538 13308 16562
rect 13308 16538 13320 16562
rect 13268 16510 13320 16538
rect 9404 16396 9456 16448
rect 10968 16396 11020 16448
rect 13084 16396 13136 16448
rect 13176 16396 13228 16448
rect 14004 16532 14056 16584
rect 15568 16668 15620 16720
rect 15108 16575 15160 16584
rect 15108 16541 15117 16575
rect 15117 16541 15151 16575
rect 15151 16541 15160 16575
rect 15108 16532 15160 16541
rect 15292 16575 15344 16584
rect 15292 16541 15301 16575
rect 15301 16541 15335 16575
rect 15335 16541 15344 16575
rect 15752 16575 15804 16584
rect 15292 16532 15344 16541
rect 15752 16541 15761 16575
rect 15761 16541 15795 16575
rect 15795 16541 15804 16575
rect 15752 16532 15804 16541
rect 17132 16600 17184 16652
rect 16856 16575 16908 16584
rect 16856 16541 16865 16575
rect 16865 16541 16899 16575
rect 16899 16541 16908 16575
rect 16856 16532 16908 16541
rect 17040 16575 17092 16584
rect 17040 16541 17054 16575
rect 17054 16541 17088 16575
rect 17088 16541 17092 16575
rect 17040 16532 17092 16541
rect 17592 16532 17644 16584
rect 18144 16668 18196 16720
rect 18144 16575 18196 16584
rect 18144 16541 18153 16575
rect 18153 16541 18187 16575
rect 18187 16541 18196 16575
rect 18144 16532 18196 16541
rect 21456 16711 21508 16720
rect 21456 16677 21465 16711
rect 21465 16677 21499 16711
rect 21499 16677 21508 16711
rect 21456 16668 21508 16677
rect 25044 16736 25096 16788
rect 29828 16736 29880 16788
rect 32496 16736 32548 16788
rect 35808 16736 35860 16788
rect 31668 16711 31720 16720
rect 20536 16532 20588 16584
rect 20628 16532 20680 16584
rect 20812 16532 20864 16584
rect 22192 16600 22244 16652
rect 21640 16575 21692 16584
rect 21640 16541 21649 16575
rect 21649 16541 21683 16575
rect 21683 16541 21692 16575
rect 21640 16532 21692 16541
rect 21732 16575 21784 16584
rect 21732 16541 21741 16575
rect 21741 16541 21775 16575
rect 21775 16541 21784 16575
rect 21732 16532 21784 16541
rect 23480 16532 23532 16584
rect 24584 16575 24636 16584
rect 22560 16464 22612 16516
rect 23296 16464 23348 16516
rect 23388 16464 23440 16516
rect 24584 16541 24593 16575
rect 24593 16541 24627 16575
rect 24627 16541 24636 16575
rect 24584 16532 24636 16541
rect 31668 16677 31677 16711
rect 31677 16677 31711 16711
rect 31711 16677 31720 16711
rect 31668 16668 31720 16677
rect 27068 16600 27120 16652
rect 27252 16643 27304 16652
rect 27252 16609 27261 16643
rect 27261 16609 27295 16643
rect 27295 16609 27304 16643
rect 27252 16600 27304 16609
rect 30472 16600 30524 16652
rect 30840 16643 30892 16652
rect 30840 16609 30849 16643
rect 30849 16609 30883 16643
rect 30883 16609 30892 16643
rect 30840 16600 30892 16609
rect 26148 16532 26200 16584
rect 29920 16575 29972 16584
rect 13452 16396 13504 16448
rect 15476 16396 15528 16448
rect 16212 16396 16264 16448
rect 16396 16396 16448 16448
rect 17040 16396 17092 16448
rect 17960 16396 18012 16448
rect 20076 16396 20128 16448
rect 23112 16396 23164 16448
rect 27620 16464 27672 16516
rect 24400 16439 24452 16448
rect 24400 16405 24409 16439
rect 24409 16405 24443 16439
rect 24443 16405 24452 16439
rect 24400 16396 24452 16405
rect 28356 16396 28408 16448
rect 29920 16541 29929 16575
rect 29929 16541 29963 16575
rect 29963 16541 29972 16575
rect 29920 16532 29972 16541
rect 30748 16575 30800 16584
rect 30748 16541 30757 16575
rect 30757 16541 30791 16575
rect 30791 16541 30800 16575
rect 30748 16532 30800 16541
rect 30932 16532 30984 16584
rect 31300 16575 31352 16584
rect 31300 16541 31309 16575
rect 31309 16541 31343 16575
rect 31343 16541 31352 16575
rect 31300 16532 31352 16541
rect 33048 16532 33100 16584
rect 33600 16600 33652 16652
rect 34796 16600 34848 16652
rect 31116 16464 31168 16516
rect 31484 16507 31536 16516
rect 31484 16473 31493 16507
rect 31493 16473 31527 16507
rect 31527 16473 31536 16507
rect 31484 16464 31536 16473
rect 31668 16464 31720 16516
rect 32128 16507 32180 16516
rect 32128 16473 32137 16507
rect 32137 16473 32171 16507
rect 32171 16473 32180 16507
rect 32128 16464 32180 16473
rect 32404 16464 32456 16516
rect 30748 16396 30800 16448
rect 31760 16396 31812 16448
rect 32864 16396 32916 16448
rect 34704 16464 34756 16516
rect 33692 16396 33744 16448
rect 34428 16396 34480 16448
rect 36544 16396 36596 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 4712 16124 4764 16176
rect 5816 16167 5868 16176
rect 5816 16133 5825 16167
rect 5825 16133 5859 16167
rect 5859 16133 5868 16167
rect 5816 16124 5868 16133
rect 7840 16192 7892 16244
rect 9128 16192 9180 16244
rect 9404 16192 9456 16244
rect 11796 16192 11848 16244
rect 15936 16192 15988 16244
rect 20168 16192 20220 16244
rect 21732 16192 21784 16244
rect 22008 16235 22060 16244
rect 22008 16201 22017 16235
rect 22017 16201 22051 16235
rect 22051 16201 22060 16235
rect 22008 16192 22060 16201
rect 2688 16099 2740 16108
rect 2688 16065 2697 16099
rect 2697 16065 2731 16099
rect 2731 16065 2740 16099
rect 2688 16056 2740 16065
rect 4804 15895 4856 15904
rect 4804 15861 4813 15895
rect 4813 15861 4847 15895
rect 4847 15861 4856 15895
rect 4804 15852 4856 15861
rect 5356 16056 5408 16108
rect 6000 16056 6052 16108
rect 6368 16099 6420 16108
rect 6368 16065 6377 16099
rect 6377 16065 6411 16099
rect 6411 16065 6420 16099
rect 6368 16056 6420 16065
rect 6276 15988 6328 16040
rect 5080 15920 5132 15972
rect 6644 15920 6696 15972
rect 8024 16124 8076 16176
rect 8208 16167 8260 16176
rect 8208 16133 8242 16167
rect 8242 16133 8260 16167
rect 8208 16124 8260 16133
rect 7380 16099 7432 16108
rect 7380 16065 7389 16099
rect 7389 16065 7423 16099
rect 7423 16065 7432 16099
rect 7380 16056 7432 16065
rect 6828 15988 6880 16040
rect 10508 15988 10560 16040
rect 10784 16099 10836 16108
rect 10784 16065 10798 16099
rect 10798 16065 10832 16099
rect 10832 16065 10836 16099
rect 12624 16124 12676 16176
rect 14924 16124 14976 16176
rect 10784 16056 10836 16065
rect 12716 16056 12768 16108
rect 17316 16124 17368 16176
rect 17868 16124 17920 16176
rect 19340 16124 19392 16176
rect 17040 16099 17092 16108
rect 17040 16065 17074 16099
rect 17074 16065 17092 16099
rect 17040 16056 17092 16065
rect 11152 15988 11204 16040
rect 6920 15852 6972 15904
rect 7288 15852 7340 15904
rect 10324 15895 10376 15904
rect 10324 15861 10333 15895
rect 10333 15861 10367 15895
rect 10367 15861 10376 15895
rect 10324 15852 10376 15861
rect 10692 15920 10744 15972
rect 13452 15920 13504 15972
rect 13544 15895 13596 15904
rect 13544 15861 13553 15895
rect 13553 15861 13587 15895
rect 13587 15861 13596 15895
rect 13544 15852 13596 15861
rect 20076 16124 20128 16176
rect 23112 16124 23164 16176
rect 23480 16192 23532 16244
rect 24676 16192 24728 16244
rect 28632 16192 28684 16244
rect 31484 16192 31536 16244
rect 23848 16124 23900 16176
rect 24400 16124 24452 16176
rect 25044 16124 25096 16176
rect 27528 16167 27580 16176
rect 27528 16133 27537 16167
rect 27537 16133 27571 16167
rect 27571 16133 27580 16167
rect 27528 16124 27580 16133
rect 30288 16124 30340 16176
rect 20628 16099 20680 16108
rect 20628 16065 20637 16099
rect 20637 16065 20671 16099
rect 20671 16065 20680 16099
rect 20628 16056 20680 16065
rect 22468 16056 22520 16108
rect 21916 15988 21968 16040
rect 26148 16056 26200 16108
rect 27068 16056 27120 16108
rect 24860 15988 24912 16040
rect 20076 15920 20128 15972
rect 20904 15920 20956 15972
rect 22468 15920 22520 15972
rect 24492 15920 24544 15972
rect 28356 16056 28408 16108
rect 28448 16056 28500 16108
rect 28908 16099 28960 16108
rect 28908 16065 28917 16099
rect 28917 16065 28951 16099
rect 28951 16065 28960 16099
rect 28908 16056 28960 16065
rect 28172 15988 28224 16040
rect 28540 15988 28592 16040
rect 30932 15988 30984 16040
rect 27896 15920 27948 15972
rect 32404 16056 32456 16108
rect 32312 15920 32364 15972
rect 15292 15852 15344 15904
rect 21088 15852 21140 15904
rect 22560 15895 22612 15904
rect 22560 15861 22569 15895
rect 22569 15861 22603 15895
rect 22603 15861 22612 15895
rect 22560 15852 22612 15861
rect 23480 15852 23532 15904
rect 27712 15852 27764 15904
rect 28172 15895 28224 15904
rect 28172 15861 28181 15895
rect 28181 15861 28215 15895
rect 28215 15861 28224 15895
rect 30748 15895 30800 15904
rect 28172 15852 28224 15861
rect 30748 15861 30757 15895
rect 30757 15861 30791 15895
rect 30791 15861 30800 15895
rect 30748 15852 30800 15861
rect 32496 15852 32548 15904
rect 34428 16056 34480 16108
rect 34612 16056 34664 16108
rect 36452 16056 36504 16108
rect 32680 16031 32732 16040
rect 32680 15997 32689 16031
rect 32689 15997 32723 16031
rect 32723 15997 32732 16031
rect 32680 15988 32732 15997
rect 33692 15920 33744 15972
rect 34244 15852 34296 15904
rect 35716 15852 35768 15904
rect 35900 15895 35952 15904
rect 35900 15861 35909 15895
rect 35909 15861 35943 15895
rect 35943 15861 35952 15895
rect 35900 15852 35952 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 1860 15555 1912 15564
rect 1860 15521 1869 15555
rect 1869 15521 1903 15555
rect 1903 15521 1912 15555
rect 1860 15512 1912 15521
rect 6736 15512 6788 15564
rect 3792 15487 3844 15496
rect 3792 15453 3801 15487
rect 3801 15453 3835 15487
rect 3835 15453 3844 15487
rect 3792 15444 3844 15453
rect 6828 15444 6880 15496
rect 3884 15376 3936 15428
rect 4804 15376 4856 15428
rect 5908 15419 5960 15428
rect 5908 15385 5942 15419
rect 5942 15385 5960 15419
rect 5908 15376 5960 15385
rect 6000 15376 6052 15428
rect 9772 15648 9824 15700
rect 10876 15648 10928 15700
rect 11152 15648 11204 15700
rect 12716 15691 12768 15700
rect 12716 15657 12725 15691
rect 12725 15657 12759 15691
rect 12759 15657 12768 15691
rect 12716 15648 12768 15657
rect 15108 15648 15160 15700
rect 15384 15648 15436 15700
rect 18144 15648 18196 15700
rect 18604 15648 18656 15700
rect 20628 15648 20680 15700
rect 23296 15691 23348 15700
rect 23296 15657 23305 15691
rect 23305 15657 23339 15691
rect 23339 15657 23348 15691
rect 23296 15648 23348 15657
rect 26148 15691 26200 15700
rect 26148 15657 26157 15691
rect 26157 15657 26191 15691
rect 26191 15657 26200 15691
rect 26148 15648 26200 15657
rect 27620 15691 27672 15700
rect 27620 15657 27629 15691
rect 27629 15657 27663 15691
rect 27663 15657 27672 15691
rect 27620 15648 27672 15657
rect 10784 15580 10836 15632
rect 11244 15580 11296 15632
rect 8944 15444 8996 15496
rect 9772 15487 9824 15496
rect 9772 15453 9781 15487
rect 9781 15453 9815 15487
rect 9815 15453 9824 15487
rect 9772 15444 9824 15453
rect 10324 15444 10376 15496
rect 10508 15444 10560 15496
rect 12072 15444 12124 15496
rect 12900 15444 12952 15496
rect 13268 15512 13320 15564
rect 14096 15512 14148 15564
rect 13176 15487 13228 15496
rect 13176 15453 13185 15487
rect 13185 15453 13219 15487
rect 13219 15453 13228 15487
rect 13176 15444 13228 15453
rect 6552 15308 6604 15360
rect 7012 15351 7064 15360
rect 7012 15317 7021 15351
rect 7021 15317 7055 15351
rect 7055 15317 7064 15351
rect 7012 15308 7064 15317
rect 11612 15419 11664 15428
rect 11612 15385 11621 15419
rect 11621 15385 11655 15419
rect 11655 15385 11664 15419
rect 11612 15376 11664 15385
rect 8852 15308 8904 15360
rect 12716 15376 12768 15428
rect 14924 15444 14976 15496
rect 16028 15444 16080 15496
rect 22468 15580 22520 15632
rect 31944 15580 31996 15632
rect 20444 15512 20496 15564
rect 17868 15487 17920 15496
rect 17868 15453 17877 15487
rect 17877 15453 17911 15487
rect 17911 15453 17920 15487
rect 17868 15444 17920 15453
rect 17960 15376 18012 15428
rect 12900 15308 12952 15360
rect 16764 15308 16816 15360
rect 21088 15487 21140 15496
rect 21088 15453 21097 15487
rect 21097 15453 21131 15487
rect 21131 15453 21140 15487
rect 21088 15444 21140 15453
rect 21272 15487 21324 15496
rect 21272 15453 21281 15487
rect 21281 15453 21315 15487
rect 21315 15453 21324 15487
rect 21272 15444 21324 15453
rect 22008 15487 22060 15496
rect 22008 15453 22017 15487
rect 22017 15453 22051 15487
rect 22051 15453 22060 15487
rect 22560 15512 22612 15564
rect 22008 15444 22060 15453
rect 23480 15487 23532 15496
rect 19708 15419 19760 15428
rect 19708 15385 19717 15419
rect 19717 15385 19751 15419
rect 19751 15385 19760 15419
rect 19708 15376 19760 15385
rect 23480 15453 23489 15487
rect 23489 15453 23523 15487
rect 23523 15453 23532 15487
rect 23480 15444 23532 15453
rect 24676 15444 24728 15496
rect 26148 15487 26200 15496
rect 26148 15453 26157 15487
rect 26157 15453 26191 15487
rect 26191 15453 26200 15487
rect 26148 15444 26200 15453
rect 27528 15444 27580 15496
rect 28172 15444 28224 15496
rect 28816 15444 28868 15496
rect 30288 15487 30340 15496
rect 30288 15453 30297 15487
rect 30297 15453 30331 15487
rect 30331 15453 30340 15487
rect 30288 15444 30340 15453
rect 30840 15512 30892 15564
rect 31852 15512 31904 15564
rect 33876 15580 33928 15632
rect 36544 15555 36596 15564
rect 36544 15521 36553 15555
rect 36553 15521 36587 15555
rect 36587 15521 36596 15555
rect 36544 15512 36596 15521
rect 30840 15376 30892 15428
rect 31852 15376 31904 15428
rect 32680 15444 32732 15496
rect 20720 15308 20772 15360
rect 22100 15308 22152 15360
rect 25044 15308 25096 15360
rect 26976 15308 27028 15360
rect 31760 15308 31812 15360
rect 32128 15308 32180 15360
rect 32864 15308 32916 15360
rect 34428 15444 34480 15496
rect 34244 15376 34296 15428
rect 35992 15376 36044 15428
rect 33784 15308 33836 15360
rect 34520 15308 34572 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 3884 15104 3936 15156
rect 2688 15011 2740 15020
rect 2688 14977 2697 15011
rect 2697 14977 2731 15011
rect 2731 14977 2740 15011
rect 2688 14968 2740 14977
rect 6000 15036 6052 15088
rect 7380 15104 7432 15156
rect 8024 15147 8076 15156
rect 8024 15113 8033 15147
rect 8033 15113 8067 15147
rect 8067 15113 8076 15147
rect 8024 15104 8076 15113
rect 8208 15104 8260 15156
rect 13268 15104 13320 15156
rect 6920 15036 6972 15088
rect 5356 14968 5408 15020
rect 5540 14968 5592 15020
rect 6368 15011 6420 15020
rect 6368 14977 6377 15011
rect 6377 14977 6411 15011
rect 6411 14977 6420 15011
rect 6368 14968 6420 14977
rect 6644 14900 6696 14952
rect 7840 14968 7892 15020
rect 8944 14968 8996 15020
rect 9036 14968 9088 15020
rect 11612 15036 11664 15088
rect 13544 15036 13596 15088
rect 11796 14968 11848 15020
rect 20996 15104 21048 15156
rect 21272 15104 21324 15156
rect 16672 15036 16724 15088
rect 7932 14900 7984 14952
rect 4804 14832 4856 14884
rect 15660 14900 15712 14952
rect 10600 14832 10652 14884
rect 17408 14900 17460 14952
rect 6460 14764 6512 14816
rect 6644 14764 6696 14816
rect 8208 14764 8260 14816
rect 15200 14764 15252 14816
rect 15476 14807 15528 14816
rect 15476 14773 15485 14807
rect 15485 14773 15519 14807
rect 15519 14773 15528 14807
rect 15476 14764 15528 14773
rect 16856 14764 16908 14816
rect 17868 14764 17920 14816
rect 18144 14900 18196 14952
rect 18328 15011 18380 15020
rect 18328 14977 18337 15011
rect 18337 14977 18371 15011
rect 18371 14977 18380 15011
rect 18328 14968 18380 14977
rect 18604 14968 18656 15020
rect 19156 14900 19208 14952
rect 20168 15036 20220 15088
rect 21272 14968 21324 15020
rect 22192 15036 22244 15088
rect 22100 15011 22152 15020
rect 22100 14977 22134 15011
rect 22134 14977 22152 15011
rect 32864 15104 32916 15156
rect 33140 15104 33192 15156
rect 33416 15104 33468 15156
rect 30472 15036 30524 15088
rect 22100 14968 22152 14977
rect 23848 15011 23900 15020
rect 19340 14900 19392 14952
rect 20536 14900 20588 14952
rect 23848 14977 23857 15011
rect 23857 14977 23891 15011
rect 23891 14977 23900 15011
rect 23848 14968 23900 14977
rect 25596 15011 25648 15020
rect 25596 14977 25605 15011
rect 25605 14977 25639 15011
rect 25639 14977 25648 15011
rect 25596 14968 25648 14977
rect 26148 14968 26200 15020
rect 28448 14968 28500 15020
rect 29000 14968 29052 15020
rect 30564 14968 30616 15020
rect 34428 14968 34480 15020
rect 32680 14943 32732 14952
rect 32680 14909 32689 14943
rect 32689 14909 32723 14943
rect 32723 14909 32732 14943
rect 32680 14900 32732 14909
rect 33968 14900 34020 14952
rect 35808 14968 35860 15020
rect 29552 14832 29604 14884
rect 19432 14764 19484 14816
rect 20168 14764 20220 14816
rect 22008 14764 22060 14816
rect 24308 14764 24360 14816
rect 26608 14764 26660 14816
rect 29644 14764 29696 14816
rect 29920 14764 29972 14816
rect 31576 14764 31628 14816
rect 31852 14764 31904 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 4712 14560 4764 14612
rect 8116 14560 8168 14612
rect 12440 14560 12492 14612
rect 14832 14560 14884 14612
rect 18328 14560 18380 14612
rect 20076 14560 20128 14612
rect 20444 14560 20496 14612
rect 20904 14560 20956 14612
rect 21916 14560 21968 14612
rect 24860 14560 24912 14612
rect 27896 14560 27948 14612
rect 5356 14492 5408 14544
rect 3792 14467 3844 14476
rect 3792 14433 3801 14467
rect 3801 14433 3835 14467
rect 3835 14433 3844 14467
rect 3792 14424 3844 14433
rect 2688 14356 2740 14408
rect 4620 14356 4672 14408
rect 6184 14424 6236 14476
rect 8208 14424 8260 14476
rect 9772 14467 9824 14476
rect 9772 14433 9781 14467
rect 9781 14433 9815 14467
rect 9815 14433 9824 14467
rect 9772 14424 9824 14433
rect 8392 14356 8444 14408
rect 9128 14399 9180 14408
rect 9128 14365 9137 14399
rect 9137 14365 9171 14399
rect 9171 14365 9180 14399
rect 9128 14356 9180 14365
rect 12072 14399 12124 14408
rect 12072 14365 12081 14399
rect 12081 14365 12115 14399
rect 12115 14365 12124 14399
rect 12072 14356 12124 14365
rect 6828 14220 6880 14272
rect 7840 14331 7892 14340
rect 7840 14297 7849 14331
rect 7849 14297 7883 14331
rect 7883 14297 7892 14331
rect 7840 14288 7892 14297
rect 11612 14288 11664 14340
rect 13176 14288 13228 14340
rect 8944 14263 8996 14272
rect 8944 14229 8953 14263
rect 8953 14229 8987 14263
rect 8987 14229 8996 14263
rect 8944 14220 8996 14229
rect 10324 14220 10376 14272
rect 15568 14492 15620 14544
rect 16488 14492 16540 14544
rect 15200 14424 15252 14476
rect 15384 14399 15436 14408
rect 15384 14365 15393 14399
rect 15393 14365 15427 14399
rect 15427 14365 15436 14399
rect 15384 14356 15436 14365
rect 16212 14424 16264 14476
rect 16672 14356 16724 14408
rect 17500 14399 17552 14408
rect 17500 14365 17509 14399
rect 17509 14365 17543 14399
rect 17543 14365 17552 14399
rect 17500 14356 17552 14365
rect 17868 14399 17920 14408
rect 17868 14365 17877 14399
rect 17877 14365 17911 14399
rect 17911 14365 17920 14399
rect 17868 14356 17920 14365
rect 15660 14288 15712 14340
rect 16856 14288 16908 14340
rect 23020 14492 23072 14544
rect 29000 14560 29052 14612
rect 34612 14560 34664 14612
rect 35900 14560 35952 14612
rect 26148 14424 26200 14476
rect 28264 14467 28316 14476
rect 28264 14433 28273 14467
rect 28273 14433 28307 14467
rect 28307 14433 28316 14467
rect 28264 14424 28316 14433
rect 19340 14356 19392 14408
rect 19432 14331 19484 14340
rect 19432 14297 19441 14331
rect 19441 14297 19475 14331
rect 19475 14297 19484 14331
rect 20076 14356 20128 14408
rect 20444 14356 20496 14408
rect 22008 14356 22060 14408
rect 22744 14356 22796 14408
rect 26976 14399 27028 14408
rect 26976 14365 26985 14399
rect 26985 14365 27019 14399
rect 27019 14365 27028 14399
rect 26976 14356 27028 14365
rect 27160 14399 27212 14408
rect 27160 14365 27169 14399
rect 27169 14365 27203 14399
rect 27203 14365 27212 14399
rect 27160 14356 27212 14365
rect 27988 14399 28040 14408
rect 27988 14365 27997 14399
rect 27997 14365 28031 14399
rect 28031 14365 28040 14399
rect 27988 14356 28040 14365
rect 29092 14424 29144 14476
rect 29552 14467 29604 14476
rect 29552 14433 29561 14467
rect 29561 14433 29595 14467
rect 29595 14433 29604 14467
rect 29552 14424 29604 14433
rect 19432 14288 19484 14297
rect 15108 14220 15160 14272
rect 17408 14220 17460 14272
rect 19340 14263 19392 14272
rect 19340 14229 19355 14263
rect 19355 14229 19389 14263
rect 19389 14229 19392 14263
rect 19340 14220 19392 14229
rect 23940 14288 23992 14340
rect 24768 14331 24820 14340
rect 24768 14297 24777 14331
rect 24777 14297 24811 14331
rect 24811 14297 24820 14331
rect 24768 14288 24820 14297
rect 27528 14288 27580 14340
rect 29644 14356 29696 14408
rect 31576 14399 31628 14408
rect 31576 14365 31585 14399
rect 31585 14365 31619 14399
rect 31619 14365 31628 14399
rect 31576 14356 31628 14365
rect 32680 14424 32732 14476
rect 34428 14424 34480 14476
rect 20904 14220 20956 14272
rect 23112 14220 23164 14272
rect 27068 14263 27120 14272
rect 27068 14229 27077 14263
rect 27077 14229 27111 14263
rect 27111 14229 27120 14263
rect 27068 14220 27120 14229
rect 28264 14263 28316 14272
rect 28264 14229 28273 14263
rect 28273 14229 28307 14263
rect 28307 14229 28316 14263
rect 28264 14220 28316 14229
rect 29552 14288 29604 14340
rect 32128 14331 32180 14340
rect 32128 14297 32137 14331
rect 32137 14297 32171 14331
rect 32171 14297 32180 14331
rect 32128 14288 32180 14297
rect 32404 14288 32456 14340
rect 32772 14288 32824 14340
rect 34520 14288 34572 14340
rect 34796 14356 34848 14408
rect 36084 14356 36136 14408
rect 32036 14220 32088 14272
rect 33324 14263 33376 14272
rect 33324 14229 33333 14263
rect 33333 14229 33367 14263
rect 33367 14229 33376 14263
rect 33324 14220 33376 14229
rect 33416 14220 33468 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 5632 14016 5684 14068
rect 6276 14016 6328 14068
rect 7104 14016 7156 14068
rect 11612 14059 11664 14068
rect 11612 14025 11621 14059
rect 11621 14025 11655 14059
rect 11655 14025 11664 14059
rect 11612 14016 11664 14025
rect 13176 14059 13228 14068
rect 13176 14025 13185 14059
rect 13185 14025 13219 14059
rect 13219 14025 13228 14059
rect 13176 14016 13228 14025
rect 15384 14016 15436 14068
rect 18052 14016 18104 14068
rect 20444 14059 20496 14068
rect 20444 14025 20453 14059
rect 20453 14025 20487 14059
rect 20487 14025 20496 14059
rect 20444 14016 20496 14025
rect 24768 14016 24820 14068
rect 4804 13948 4856 14000
rect 2688 13923 2740 13932
rect 2688 13889 2697 13923
rect 2697 13889 2731 13923
rect 2731 13889 2740 13923
rect 2688 13880 2740 13889
rect 6644 13948 6696 14000
rect 7012 13948 7064 14000
rect 8116 13948 8168 14000
rect 10048 13948 10100 14000
rect 12164 13948 12216 14000
rect 6368 13923 6420 13932
rect 6368 13889 6377 13923
rect 6377 13889 6411 13923
rect 6411 13889 6420 13923
rect 6368 13880 6420 13889
rect 6552 13923 6604 13932
rect 6552 13889 6561 13923
rect 6561 13889 6595 13923
rect 6595 13889 6604 13923
rect 6552 13880 6604 13889
rect 7196 13923 7248 13932
rect 7196 13889 7205 13923
rect 7205 13889 7239 13923
rect 7239 13889 7248 13923
rect 7196 13880 7248 13889
rect 7840 13880 7892 13932
rect 8208 13923 8260 13932
rect 8208 13889 8217 13923
rect 8217 13889 8251 13923
rect 8251 13889 8260 13923
rect 8208 13880 8260 13889
rect 8300 13880 8352 13932
rect 5724 13812 5776 13864
rect 6736 13812 6788 13864
rect 9220 13923 9272 13932
rect 9220 13889 9229 13923
rect 9229 13889 9263 13923
rect 9263 13889 9272 13923
rect 9220 13880 9272 13889
rect 10508 13923 10560 13932
rect 10508 13889 10517 13923
rect 10517 13889 10551 13923
rect 10551 13889 10560 13923
rect 10508 13880 10560 13889
rect 9772 13812 9824 13864
rect 10324 13855 10376 13864
rect 10324 13821 10333 13855
rect 10333 13821 10367 13855
rect 10367 13821 10376 13855
rect 10324 13812 10376 13821
rect 11796 13880 11848 13932
rect 13268 13923 13320 13932
rect 12440 13855 12492 13864
rect 12440 13821 12449 13855
rect 12449 13821 12483 13855
rect 12483 13821 12492 13855
rect 12440 13812 12492 13821
rect 12164 13744 12216 13796
rect 13268 13889 13277 13923
rect 13277 13889 13311 13923
rect 13311 13889 13320 13923
rect 13268 13880 13320 13889
rect 15660 13948 15712 14000
rect 17316 13948 17368 14000
rect 19340 13991 19392 14000
rect 15108 13923 15160 13932
rect 15108 13889 15117 13923
rect 15117 13889 15151 13923
rect 15151 13889 15160 13923
rect 15108 13880 15160 13889
rect 15476 13923 15528 13932
rect 15476 13889 15485 13923
rect 15485 13889 15519 13923
rect 15519 13889 15528 13923
rect 15476 13880 15528 13889
rect 15844 13923 15896 13932
rect 15844 13889 15853 13923
rect 15853 13889 15887 13923
rect 15887 13889 15896 13923
rect 15844 13880 15896 13889
rect 13176 13744 13228 13796
rect 15568 13812 15620 13864
rect 17224 13880 17276 13932
rect 19340 13957 19374 13991
rect 19374 13957 19392 13991
rect 19340 13948 19392 13957
rect 21548 13880 21600 13932
rect 22744 13948 22796 14000
rect 22192 13880 22244 13932
rect 23664 13880 23716 13932
rect 24860 13948 24912 14000
rect 25596 13948 25648 14000
rect 27068 13880 27120 13932
rect 27712 13880 27764 13932
rect 27988 13880 28040 13932
rect 17500 13812 17552 13864
rect 17776 13812 17828 13864
rect 17868 13855 17920 13864
rect 17868 13821 17877 13855
rect 17877 13821 17911 13855
rect 17911 13821 17920 13855
rect 17868 13812 17920 13821
rect 20168 13812 20220 13864
rect 20352 13812 20404 13864
rect 15108 13744 15160 13796
rect 17960 13787 18012 13796
rect 17960 13753 17969 13787
rect 17969 13753 18003 13787
rect 18003 13753 18012 13787
rect 17960 13744 18012 13753
rect 10416 13719 10468 13728
rect 10416 13685 10425 13719
rect 10425 13685 10459 13719
rect 10459 13685 10468 13719
rect 10416 13676 10468 13685
rect 15476 13676 15528 13728
rect 24400 13676 24452 13728
rect 26056 13676 26108 13728
rect 26240 13676 26292 13728
rect 30656 14016 30708 14068
rect 32864 14016 32916 14068
rect 34244 14016 34296 14068
rect 35716 14016 35768 14068
rect 30840 13948 30892 14000
rect 32588 13948 32640 14000
rect 29092 13923 29144 13932
rect 29092 13889 29101 13923
rect 29101 13889 29135 13923
rect 29135 13889 29144 13923
rect 29092 13880 29144 13889
rect 29920 13923 29972 13932
rect 29920 13889 29929 13923
rect 29929 13889 29963 13923
rect 29963 13889 29972 13923
rect 29920 13880 29972 13889
rect 30748 13880 30800 13932
rect 31668 13880 31720 13932
rect 32680 13880 32732 13932
rect 33140 13923 33192 13932
rect 33140 13889 33149 13923
rect 33149 13889 33183 13923
rect 33183 13889 33192 13923
rect 33140 13880 33192 13889
rect 34428 13880 34480 13932
rect 34612 13880 34664 13932
rect 34152 13812 34204 13864
rect 34704 13676 34756 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 5448 13472 5500 13524
rect 9128 13472 9180 13524
rect 9220 13404 9272 13456
rect 6460 13311 6512 13320
rect 6460 13277 6469 13311
rect 6469 13277 6503 13311
rect 6503 13277 6512 13311
rect 6460 13268 6512 13277
rect 6828 13268 6880 13320
rect 7932 13200 7984 13252
rect 8852 13200 8904 13252
rect 9128 13243 9180 13252
rect 9128 13209 9137 13243
rect 9137 13209 9171 13243
rect 9171 13209 9180 13243
rect 9128 13200 9180 13209
rect 10324 13243 10376 13252
rect 10324 13209 10358 13243
rect 10358 13209 10376 13243
rect 10324 13200 10376 13209
rect 10232 13132 10284 13184
rect 13636 13472 13688 13524
rect 15200 13472 15252 13524
rect 14464 13404 14516 13456
rect 16948 13472 17000 13524
rect 23664 13515 23716 13524
rect 16672 13404 16724 13456
rect 17868 13404 17920 13456
rect 12072 13379 12124 13388
rect 12072 13345 12081 13379
rect 12081 13345 12115 13379
rect 12115 13345 12124 13379
rect 12072 13336 12124 13345
rect 14004 13336 14056 13388
rect 12900 13200 12952 13252
rect 14096 13311 14148 13320
rect 14096 13277 14105 13311
rect 14105 13277 14139 13311
rect 14139 13277 14148 13311
rect 17408 13336 17460 13388
rect 19340 13404 19392 13456
rect 23664 13481 23673 13515
rect 23673 13481 23707 13515
rect 23707 13481 23716 13515
rect 23664 13472 23716 13481
rect 24492 13515 24544 13524
rect 24492 13481 24501 13515
rect 24501 13481 24535 13515
rect 24535 13481 24544 13515
rect 26424 13515 26476 13524
rect 24492 13472 24544 13481
rect 21548 13404 21600 13456
rect 14096 13268 14148 13277
rect 15108 13268 15160 13320
rect 15476 13311 15528 13320
rect 15476 13277 15485 13311
rect 15485 13277 15519 13311
rect 15519 13277 15528 13311
rect 15476 13268 15528 13277
rect 15568 13311 15620 13320
rect 15568 13277 15577 13311
rect 15577 13277 15611 13311
rect 15611 13277 15620 13311
rect 15936 13311 15988 13320
rect 15568 13268 15620 13277
rect 15936 13277 15945 13311
rect 15945 13277 15979 13311
rect 15979 13277 15988 13311
rect 15936 13268 15988 13277
rect 16764 13268 16816 13320
rect 17132 13311 17184 13320
rect 17132 13277 17138 13311
rect 17138 13277 17184 13311
rect 17132 13268 17184 13277
rect 17868 13268 17920 13320
rect 15292 13200 15344 13252
rect 16120 13200 16172 13252
rect 18788 13200 18840 13252
rect 20536 13336 20588 13388
rect 19432 13311 19484 13320
rect 19432 13277 19441 13311
rect 19441 13277 19475 13311
rect 19475 13277 19484 13311
rect 19432 13268 19484 13277
rect 24400 13311 24452 13320
rect 19156 13200 19208 13252
rect 23756 13200 23808 13252
rect 24400 13277 24409 13311
rect 24409 13277 24443 13311
rect 24443 13277 24452 13311
rect 24400 13268 24452 13277
rect 24952 13336 25004 13388
rect 26424 13481 26433 13515
rect 26433 13481 26467 13515
rect 26467 13481 26476 13515
rect 26424 13472 26476 13481
rect 27160 13472 27212 13524
rect 27712 13515 27764 13524
rect 27712 13481 27721 13515
rect 27721 13481 27755 13515
rect 27755 13481 27764 13515
rect 27712 13472 27764 13481
rect 31668 13472 31720 13524
rect 34612 13472 34664 13524
rect 26056 13404 26108 13456
rect 26516 13379 26568 13388
rect 25044 13268 25096 13320
rect 26240 13311 26292 13320
rect 26240 13277 26249 13311
rect 26249 13277 26283 13311
rect 26283 13277 26292 13311
rect 26240 13268 26292 13277
rect 26516 13345 26525 13379
rect 26525 13345 26559 13379
rect 26559 13345 26568 13379
rect 26516 13336 26568 13345
rect 27252 13379 27304 13388
rect 27252 13345 27261 13379
rect 27261 13345 27295 13379
rect 27295 13345 27304 13379
rect 27252 13336 27304 13345
rect 26976 13311 27028 13320
rect 26976 13277 26985 13311
rect 26985 13277 27019 13311
rect 27019 13277 27028 13311
rect 26976 13268 27028 13277
rect 27528 13268 27580 13320
rect 28264 13268 28316 13320
rect 30472 13311 30524 13320
rect 30472 13277 30481 13311
rect 30481 13277 30515 13311
rect 30515 13277 30524 13311
rect 30472 13268 30524 13277
rect 35992 13472 36044 13524
rect 31852 13268 31904 13320
rect 33324 13268 33376 13320
rect 33600 13311 33652 13320
rect 33600 13277 33609 13311
rect 33609 13277 33643 13311
rect 33643 13277 33652 13311
rect 33600 13268 33652 13277
rect 34152 13268 34204 13320
rect 26884 13200 26936 13252
rect 32864 13200 32916 13252
rect 19432 13132 19484 13184
rect 25688 13175 25740 13184
rect 25688 13141 25697 13175
rect 25697 13141 25731 13175
rect 25731 13141 25740 13175
rect 25688 13132 25740 13141
rect 30288 13175 30340 13184
rect 30288 13141 30297 13175
rect 30297 13141 30331 13175
rect 30331 13141 30340 13175
rect 30288 13132 30340 13141
rect 32772 13132 32824 13184
rect 33692 13132 33744 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 6092 12928 6144 12980
rect 8392 12928 8444 12980
rect 9036 12928 9088 12980
rect 3700 12860 3752 12912
rect 8944 12860 8996 12912
rect 12900 12903 12952 12912
rect 12900 12869 12909 12903
rect 12909 12869 12943 12903
rect 12943 12869 12952 12903
rect 12900 12860 12952 12869
rect 14096 12860 14148 12912
rect 16396 12860 16448 12912
rect 17040 12860 17092 12912
rect 17592 12860 17644 12912
rect 17684 12860 17736 12912
rect 19340 12903 19392 12912
rect 19340 12869 19349 12903
rect 19349 12869 19383 12903
rect 19383 12869 19392 12903
rect 19984 12903 20036 12912
rect 19340 12860 19392 12869
rect 19984 12869 19993 12903
rect 19993 12869 20027 12903
rect 20027 12869 20036 12903
rect 19984 12860 20036 12869
rect 2688 12835 2740 12844
rect 2688 12801 2697 12835
rect 2697 12801 2731 12835
rect 2731 12801 2740 12835
rect 2688 12792 2740 12801
rect 6828 12792 6880 12844
rect 5264 12724 5316 12776
rect 12808 12835 12860 12844
rect 12808 12801 12817 12835
rect 12817 12801 12851 12835
rect 12851 12801 12860 12835
rect 12808 12792 12860 12801
rect 10048 12767 10100 12776
rect 10048 12733 10057 12767
rect 10057 12733 10091 12767
rect 10091 12733 10100 12767
rect 10048 12724 10100 12733
rect 10232 12767 10284 12776
rect 10232 12733 10241 12767
rect 10241 12733 10275 12767
rect 10275 12733 10284 12767
rect 10232 12724 10284 12733
rect 10692 12724 10744 12776
rect 11796 12767 11848 12776
rect 9128 12656 9180 12708
rect 10416 12656 10468 12708
rect 10876 12656 10928 12708
rect 10232 12631 10284 12640
rect 10232 12597 10241 12631
rect 10241 12597 10275 12631
rect 10275 12597 10284 12631
rect 10232 12588 10284 12597
rect 11796 12733 11805 12767
rect 11805 12733 11839 12767
rect 11839 12733 11848 12767
rect 11796 12724 11848 12733
rect 13268 12792 13320 12844
rect 14004 12792 14056 12844
rect 15200 12835 15252 12844
rect 15200 12801 15209 12835
rect 15209 12801 15243 12835
rect 15243 12801 15252 12835
rect 15200 12792 15252 12801
rect 16672 12835 16724 12844
rect 16672 12801 16681 12835
rect 16681 12801 16715 12835
rect 16715 12801 16724 12835
rect 16672 12792 16724 12801
rect 15936 12656 15988 12708
rect 16396 12724 16448 12776
rect 18052 12835 18104 12844
rect 18052 12801 18061 12835
rect 18061 12801 18095 12835
rect 18095 12801 18104 12835
rect 18052 12792 18104 12801
rect 18328 12792 18380 12844
rect 18604 12792 18656 12844
rect 18880 12792 18932 12844
rect 19156 12835 19208 12844
rect 19156 12801 19165 12835
rect 19165 12801 19199 12835
rect 19199 12801 19208 12835
rect 19156 12792 19208 12801
rect 19432 12835 19484 12844
rect 19432 12801 19441 12835
rect 19441 12801 19475 12835
rect 19475 12801 19484 12835
rect 19432 12792 19484 12801
rect 20536 12792 20588 12844
rect 21272 12792 21324 12844
rect 16764 12699 16816 12708
rect 15660 12588 15712 12640
rect 16396 12588 16448 12640
rect 16764 12665 16773 12699
rect 16773 12665 16807 12699
rect 16807 12665 16816 12699
rect 16764 12656 16816 12665
rect 19432 12656 19484 12708
rect 20904 12656 20956 12708
rect 20720 12631 20772 12640
rect 20720 12597 20729 12631
rect 20729 12597 20763 12631
rect 20763 12597 20772 12631
rect 20720 12588 20772 12597
rect 30288 12860 30340 12912
rect 31668 12860 31720 12912
rect 23756 12792 23808 12844
rect 25136 12792 25188 12844
rect 28264 12835 28316 12844
rect 28264 12801 28273 12835
rect 28273 12801 28307 12835
rect 28307 12801 28316 12835
rect 28264 12792 28316 12801
rect 28448 12835 28500 12844
rect 28448 12801 28457 12835
rect 28457 12801 28491 12835
rect 28491 12801 28500 12835
rect 28448 12792 28500 12801
rect 28908 12835 28960 12844
rect 28908 12801 28917 12835
rect 28917 12801 28951 12835
rect 28951 12801 28960 12835
rect 28908 12792 28960 12801
rect 28356 12724 28408 12776
rect 34060 12792 34112 12844
rect 29644 12724 29696 12776
rect 29920 12767 29972 12776
rect 29920 12733 29929 12767
rect 29929 12733 29963 12767
rect 29963 12733 29972 12767
rect 29920 12724 29972 12733
rect 29092 12656 29144 12708
rect 23480 12588 23532 12640
rect 23664 12631 23716 12640
rect 23664 12597 23673 12631
rect 23673 12597 23707 12631
rect 23707 12597 23716 12631
rect 23664 12588 23716 12597
rect 28172 12588 28224 12640
rect 28724 12588 28776 12640
rect 31300 12631 31352 12640
rect 31300 12597 31309 12631
rect 31309 12597 31343 12631
rect 31343 12597 31352 12631
rect 31300 12588 31352 12597
rect 31760 12588 31812 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 8300 12384 8352 12436
rect 10324 12427 10376 12436
rect 10324 12393 10333 12427
rect 10333 12393 10367 12427
rect 10367 12393 10376 12427
rect 10324 12384 10376 12393
rect 14280 12427 14332 12436
rect 14280 12393 14289 12427
rect 14289 12393 14323 12427
rect 14323 12393 14332 12427
rect 14280 12384 14332 12393
rect 15752 12384 15804 12436
rect 16396 12384 16448 12436
rect 16764 12384 16816 12436
rect 6828 12248 6880 12300
rect 14464 12316 14516 12368
rect 16856 12316 16908 12368
rect 17684 12384 17736 12436
rect 19800 12427 19852 12436
rect 19800 12393 19809 12427
rect 19809 12393 19843 12427
rect 19843 12393 19852 12427
rect 19800 12384 19852 12393
rect 15476 12248 15528 12300
rect 16488 12248 16540 12300
rect 17868 12316 17920 12368
rect 23480 12384 23532 12436
rect 26976 12427 27028 12436
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 10416 12223 10468 12232
rect 10416 12189 10425 12223
rect 10425 12189 10459 12223
rect 10459 12189 10468 12223
rect 10416 12180 10468 12189
rect 11796 12180 11848 12232
rect 15108 12180 15160 12232
rect 16028 12180 16080 12232
rect 17960 12180 18012 12232
rect 19248 12180 19300 12232
rect 21824 12180 21876 12232
rect 12164 12112 12216 12164
rect 14096 12155 14148 12164
rect 14096 12121 14105 12155
rect 14105 12121 14139 12155
rect 14139 12121 14148 12155
rect 14096 12112 14148 12121
rect 15384 12112 15436 12164
rect 16396 12112 16448 12164
rect 18328 12112 18380 12164
rect 20720 12155 20772 12164
rect 20720 12121 20754 12155
rect 20754 12121 20772 12155
rect 22744 12155 22796 12164
rect 20720 12112 20772 12121
rect 22744 12121 22753 12155
rect 22753 12121 22787 12155
rect 22787 12121 22796 12155
rect 22744 12112 22796 12121
rect 23020 12291 23072 12300
rect 23020 12257 23029 12291
rect 23029 12257 23063 12291
rect 23063 12257 23072 12291
rect 23020 12248 23072 12257
rect 23480 12180 23532 12232
rect 26976 12393 26985 12427
rect 26985 12393 27019 12427
rect 27019 12393 27028 12427
rect 26976 12384 27028 12393
rect 30472 12384 30524 12436
rect 32588 12384 32640 12436
rect 34152 12384 34204 12436
rect 35532 12316 35584 12368
rect 28356 12248 28408 12300
rect 24124 12180 24176 12232
rect 25136 12223 25188 12232
rect 24860 12112 24912 12164
rect 25136 12189 25145 12223
rect 25145 12189 25179 12223
rect 25179 12189 25188 12223
rect 25136 12180 25188 12189
rect 25596 12223 25648 12232
rect 25596 12189 25605 12223
rect 25605 12189 25639 12223
rect 25639 12189 25648 12223
rect 25596 12180 25648 12189
rect 25688 12180 25740 12232
rect 27804 12223 27856 12232
rect 27804 12189 27813 12223
rect 27813 12189 27847 12223
rect 27847 12189 27856 12223
rect 27804 12180 27856 12189
rect 28448 12180 28500 12232
rect 28816 12223 28868 12232
rect 28816 12189 28825 12223
rect 28825 12189 28859 12223
rect 28859 12189 28868 12223
rect 28816 12180 28868 12189
rect 32772 12248 32824 12300
rect 29552 12223 29604 12232
rect 29552 12189 29561 12223
rect 29561 12189 29595 12223
rect 29595 12189 29604 12223
rect 29552 12180 29604 12189
rect 29644 12180 29696 12232
rect 31300 12180 31352 12232
rect 26424 12112 26476 12164
rect 31852 12180 31904 12232
rect 18972 12044 19024 12096
rect 20076 12044 20128 12096
rect 24032 12044 24084 12096
rect 25964 12044 26016 12096
rect 30748 12044 30800 12096
rect 32128 12112 32180 12164
rect 33232 12112 33284 12164
rect 33600 12155 33652 12164
rect 33600 12121 33609 12155
rect 33609 12121 33643 12155
rect 33643 12121 33652 12155
rect 33600 12112 33652 12121
rect 33692 12044 33744 12096
rect 33784 12087 33836 12096
rect 33784 12053 33793 12087
rect 33793 12053 33827 12087
rect 33827 12053 33836 12087
rect 33784 12044 33836 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 7932 11883 7984 11892
rect 7932 11849 7941 11883
rect 7941 11849 7975 11883
rect 7975 11849 7984 11883
rect 7932 11840 7984 11849
rect 10876 11840 10928 11892
rect 17132 11840 17184 11892
rect 18052 11840 18104 11892
rect 19984 11840 20036 11892
rect 21364 11840 21416 11892
rect 24860 11840 24912 11892
rect 25228 11840 25280 11892
rect 28448 11840 28500 11892
rect 28724 11840 28776 11892
rect 34060 11883 34112 11892
rect 34060 11849 34069 11883
rect 34069 11849 34103 11883
rect 34103 11849 34112 11883
rect 34060 11840 34112 11849
rect 9220 11772 9272 11824
rect 16856 11815 16908 11824
rect 16856 11781 16865 11815
rect 16865 11781 16899 11815
rect 16899 11781 16908 11815
rect 16856 11772 16908 11781
rect 20536 11772 20588 11824
rect 24032 11815 24084 11824
rect 8116 11747 8168 11756
rect 8116 11713 8125 11747
rect 8125 11713 8159 11747
rect 8159 11713 8168 11747
rect 8116 11704 8168 11713
rect 12624 11747 12676 11756
rect 12624 11713 12633 11747
rect 12633 11713 12667 11747
rect 12667 11713 12676 11747
rect 12624 11704 12676 11713
rect 13544 11704 13596 11756
rect 16764 11704 16816 11756
rect 18328 11704 18380 11756
rect 18972 11704 19024 11756
rect 21088 11747 21140 11756
rect 21088 11713 21097 11747
rect 21097 11713 21131 11747
rect 21131 11713 21140 11747
rect 21088 11704 21140 11713
rect 21272 11747 21324 11756
rect 21272 11713 21281 11747
rect 21281 11713 21315 11747
rect 21315 11713 21324 11747
rect 21272 11704 21324 11713
rect 21824 11747 21876 11756
rect 21824 11713 21833 11747
rect 21833 11713 21867 11747
rect 21867 11713 21876 11747
rect 21824 11704 21876 11713
rect 24032 11781 24066 11815
rect 24066 11781 24084 11815
rect 24032 11772 24084 11781
rect 24124 11772 24176 11824
rect 12900 11679 12952 11688
rect 12900 11645 12909 11679
rect 12909 11645 12943 11679
rect 12943 11645 12952 11679
rect 12900 11636 12952 11645
rect 16120 11679 16172 11688
rect 16120 11645 16129 11679
rect 16129 11645 16163 11679
rect 16163 11645 16172 11679
rect 16120 11636 16172 11645
rect 16396 11636 16448 11688
rect 20076 11636 20128 11688
rect 24952 11704 25004 11756
rect 27620 11772 27672 11824
rect 26884 11704 26936 11756
rect 28356 11747 28408 11756
rect 25136 11636 25188 11688
rect 28356 11713 28365 11747
rect 28365 11713 28399 11747
rect 28399 11713 28408 11747
rect 28356 11704 28408 11713
rect 31760 11704 31812 11756
rect 27804 11636 27856 11688
rect 28724 11679 28776 11688
rect 28724 11645 28733 11679
rect 28733 11645 28767 11679
rect 28767 11645 28776 11679
rect 28724 11636 28776 11645
rect 33692 11704 33744 11756
rect 15752 11568 15804 11620
rect 12348 11500 12400 11552
rect 12716 11500 12768 11552
rect 13452 11500 13504 11552
rect 16488 11500 16540 11552
rect 18236 11500 18288 11552
rect 18512 11500 18564 11552
rect 19432 11568 19484 11620
rect 19708 11568 19760 11620
rect 19984 11568 20036 11620
rect 21456 11568 21508 11620
rect 32588 11636 32640 11688
rect 25688 11543 25740 11552
rect 25688 11509 25697 11543
rect 25697 11509 25731 11543
rect 25731 11509 25740 11543
rect 25688 11500 25740 11509
rect 27344 11500 27396 11552
rect 33324 11500 33376 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 15844 11296 15896 11348
rect 13452 11271 13504 11280
rect 13452 11237 13461 11271
rect 13461 11237 13495 11271
rect 13495 11237 13504 11271
rect 13452 11228 13504 11237
rect 16856 11228 16908 11280
rect 15568 11160 15620 11212
rect 15660 11160 15712 11212
rect 18328 11296 18380 11348
rect 20260 11296 20312 11348
rect 21088 11296 21140 11348
rect 21456 11339 21508 11348
rect 21456 11305 21465 11339
rect 21465 11305 21499 11339
rect 21499 11305 21508 11339
rect 21456 11296 21508 11305
rect 23020 11296 23072 11348
rect 25504 11296 25556 11348
rect 27896 11296 27948 11348
rect 10416 11092 10468 11144
rect 11520 11092 11572 11144
rect 12348 11135 12400 11144
rect 12348 11101 12382 11135
rect 12382 11101 12400 11135
rect 12348 11092 12400 11101
rect 14280 11092 14332 11144
rect 15292 11092 15344 11144
rect 18236 11228 18288 11280
rect 21916 11228 21968 11280
rect 18144 11160 18196 11212
rect 18604 11160 18656 11212
rect 23480 11228 23532 11280
rect 24400 11228 24452 11280
rect 24124 11160 24176 11212
rect 29920 11160 29972 11212
rect 32588 11228 32640 11280
rect 19248 11135 19300 11144
rect 19248 11101 19257 11135
rect 19257 11101 19291 11135
rect 19291 11101 19300 11135
rect 19248 11092 19300 11101
rect 19800 11092 19852 11144
rect 21088 11092 21140 11144
rect 21364 11092 21416 11144
rect 10784 11024 10836 11076
rect 13820 11024 13872 11076
rect 15200 11067 15252 11076
rect 15200 11033 15209 11067
rect 15209 11033 15243 11067
rect 15243 11033 15252 11067
rect 15200 11024 15252 11033
rect 15568 11024 15620 11076
rect 10048 10999 10100 11008
rect 10048 10965 10057 10999
rect 10057 10965 10091 10999
rect 10091 10965 10100 10999
rect 10048 10956 10100 10965
rect 16028 11067 16080 11076
rect 16028 11033 16037 11067
rect 16037 11033 16071 11067
rect 16071 11033 16080 11067
rect 16028 11024 16080 11033
rect 20076 11024 20128 11076
rect 20536 11024 20588 11076
rect 19340 10956 19392 11008
rect 20260 10956 20312 11008
rect 23020 11135 23072 11144
rect 23020 11101 23029 11135
rect 23029 11101 23063 11135
rect 23063 11101 23072 11135
rect 23020 11092 23072 11101
rect 25596 11092 25648 11144
rect 26240 11092 26292 11144
rect 32404 11135 32456 11144
rect 32404 11101 32413 11135
rect 32413 11101 32447 11135
rect 32447 11101 32456 11135
rect 32404 11092 32456 11101
rect 34704 11092 34756 11144
rect 25688 11024 25740 11076
rect 27528 11024 27580 11076
rect 30932 11024 30984 11076
rect 30380 10956 30432 11008
rect 30840 10956 30892 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 7564 10752 7616 10804
rect 10324 10752 10376 10804
rect 16396 10752 16448 10804
rect 16672 10752 16724 10804
rect 17224 10752 17276 10804
rect 20076 10795 20128 10804
rect 10048 10616 10100 10668
rect 10324 10616 10376 10668
rect 15016 10684 15068 10736
rect 18880 10684 18932 10736
rect 19432 10684 19484 10736
rect 20076 10761 20085 10795
rect 20085 10761 20119 10795
rect 20119 10761 20128 10795
rect 20076 10752 20128 10761
rect 21088 10752 21140 10804
rect 11520 10659 11572 10668
rect 11520 10625 11529 10659
rect 11529 10625 11563 10659
rect 11563 10625 11572 10659
rect 11520 10616 11572 10625
rect 11612 10616 11664 10668
rect 14004 10659 14056 10668
rect 14004 10625 14013 10659
rect 14013 10625 14047 10659
rect 14047 10625 14056 10659
rect 14004 10616 14056 10625
rect 11428 10548 11480 10600
rect 14280 10591 14332 10600
rect 14280 10557 14289 10591
rect 14289 10557 14323 10591
rect 14323 10557 14332 10591
rect 14280 10548 14332 10557
rect 10600 10523 10652 10532
rect 10600 10489 10609 10523
rect 10609 10489 10643 10523
rect 10643 10489 10652 10523
rect 10600 10480 10652 10489
rect 10876 10523 10928 10532
rect 10876 10489 10885 10523
rect 10885 10489 10919 10523
rect 10919 10489 10928 10523
rect 10876 10480 10928 10489
rect 12900 10523 12952 10532
rect 12900 10489 12909 10523
rect 12909 10489 12943 10523
rect 12943 10489 12952 10523
rect 15292 10616 15344 10668
rect 15660 10616 15712 10668
rect 16212 10616 16264 10668
rect 15200 10548 15252 10600
rect 16764 10659 16816 10668
rect 16764 10625 16773 10659
rect 16773 10625 16807 10659
rect 16807 10625 16816 10659
rect 16764 10616 16816 10625
rect 12900 10480 12952 10489
rect 10784 10455 10836 10464
rect 10784 10421 10793 10455
rect 10793 10421 10827 10455
rect 10827 10421 10836 10455
rect 10784 10412 10836 10421
rect 13820 10412 13872 10464
rect 16396 10412 16448 10464
rect 17592 10616 17644 10668
rect 19340 10591 19392 10600
rect 19340 10557 19349 10591
rect 19349 10557 19383 10591
rect 19383 10557 19392 10591
rect 19340 10548 19392 10557
rect 21272 10616 21324 10668
rect 21916 10616 21968 10668
rect 22744 10684 22796 10736
rect 27620 10752 27672 10804
rect 27804 10684 27856 10736
rect 25320 10616 25372 10668
rect 25504 10548 25556 10600
rect 31024 10752 31076 10804
rect 33232 10752 33284 10804
rect 29552 10684 29604 10736
rect 30472 10684 30524 10736
rect 29368 10616 29420 10668
rect 30564 10616 30616 10668
rect 32772 10684 32824 10736
rect 33324 10684 33376 10736
rect 30840 10591 30892 10600
rect 30840 10557 30849 10591
rect 30849 10557 30883 10591
rect 30883 10557 30892 10591
rect 30840 10548 30892 10557
rect 32588 10548 32640 10600
rect 26976 10480 27028 10532
rect 30380 10480 30432 10532
rect 19984 10412 20036 10464
rect 24952 10455 25004 10464
rect 24952 10421 24961 10455
rect 24961 10421 24995 10455
rect 24995 10421 25004 10455
rect 24952 10412 25004 10421
rect 25320 10412 25372 10464
rect 25596 10412 25648 10464
rect 26700 10412 26752 10464
rect 27436 10412 27488 10464
rect 28816 10412 28868 10464
rect 29552 10455 29604 10464
rect 29552 10421 29561 10455
rect 29561 10421 29595 10455
rect 29595 10421 29604 10455
rect 29552 10412 29604 10421
rect 31116 10412 31168 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 11612 10208 11664 10260
rect 14280 10208 14332 10260
rect 15200 10208 15252 10260
rect 16488 10251 16540 10260
rect 16488 10217 16497 10251
rect 16497 10217 16531 10251
rect 16531 10217 16540 10251
rect 16488 10208 16540 10217
rect 17960 10208 18012 10260
rect 18696 10208 18748 10260
rect 25872 10208 25924 10260
rect 27528 10251 27580 10260
rect 27528 10217 27537 10251
rect 27537 10217 27571 10251
rect 27571 10217 27580 10251
rect 27528 10208 27580 10217
rect 30932 10251 30984 10260
rect 30932 10217 30941 10251
rect 30941 10217 30975 10251
rect 30975 10217 30984 10251
rect 30932 10208 30984 10217
rect 33600 10208 33652 10260
rect 10600 10140 10652 10192
rect 14096 10140 14148 10192
rect 17224 10140 17276 10192
rect 26700 10140 26752 10192
rect 10692 10072 10744 10124
rect 9128 10047 9180 10056
rect 9128 10013 9137 10047
rect 9137 10013 9171 10047
rect 9171 10013 9180 10047
rect 9128 10004 9180 10013
rect 10876 10004 10928 10056
rect 11336 10004 11388 10056
rect 12716 10004 12768 10056
rect 12900 10072 12952 10124
rect 14004 10072 14056 10124
rect 32680 10140 32732 10192
rect 13820 10004 13872 10056
rect 30380 10072 30432 10124
rect 16120 10004 16172 10056
rect 19340 10004 19392 10056
rect 21916 10004 21968 10056
rect 23020 10004 23072 10056
rect 26240 10004 26292 10056
rect 27436 10047 27488 10056
rect 27436 10013 27445 10047
rect 27445 10013 27479 10047
rect 27479 10013 27488 10047
rect 27436 10004 27488 10013
rect 28816 10047 28868 10056
rect 1400 9868 1452 9920
rect 8944 9911 8996 9920
rect 8944 9877 8953 9911
rect 8953 9877 8987 9911
rect 8987 9877 8996 9911
rect 8944 9868 8996 9877
rect 9036 9868 9088 9920
rect 11244 9868 11296 9920
rect 15200 9936 15252 9988
rect 16028 9936 16080 9988
rect 16396 9979 16448 9988
rect 15016 9868 15068 9920
rect 16396 9945 16405 9979
rect 16405 9945 16439 9979
rect 16439 9945 16448 9979
rect 16396 9936 16448 9945
rect 17500 9979 17552 9988
rect 17500 9945 17534 9979
rect 17534 9945 17552 9979
rect 17500 9936 17552 9945
rect 20904 9936 20956 9988
rect 26148 9936 26200 9988
rect 28816 10013 28825 10047
rect 28825 10013 28859 10047
rect 28859 10013 28868 10047
rect 28816 10004 28868 10013
rect 30472 10004 30524 10056
rect 32036 10004 32088 10056
rect 32588 10004 32640 10056
rect 33784 10004 33836 10056
rect 16764 9868 16816 9920
rect 20720 9868 20772 9920
rect 21732 9868 21784 9920
rect 26332 9868 26384 9920
rect 28908 9911 28960 9920
rect 28908 9877 28917 9911
rect 28917 9877 28951 9911
rect 28951 9877 28960 9911
rect 28908 9868 28960 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 17500 9707 17552 9716
rect 17500 9673 17509 9707
rect 17509 9673 17543 9707
rect 17543 9673 17552 9707
rect 17500 9664 17552 9673
rect 20904 9707 20956 9716
rect 20904 9673 20913 9707
rect 20913 9673 20947 9707
rect 20947 9673 20956 9707
rect 20904 9664 20956 9673
rect 8944 9596 8996 9648
rect 12440 9596 12492 9648
rect 11060 9528 11112 9580
rect 11980 9571 12032 9580
rect 11980 9537 11989 9571
rect 11989 9537 12023 9571
rect 12023 9537 12032 9571
rect 11980 9528 12032 9537
rect 12624 9528 12676 9580
rect 7932 9503 7984 9512
rect 7932 9469 7941 9503
rect 7941 9469 7975 9503
rect 7975 9469 7984 9503
rect 7932 9460 7984 9469
rect 12716 9460 12768 9512
rect 13544 9528 13596 9580
rect 15752 9596 15804 9648
rect 20168 9596 20220 9648
rect 20628 9596 20680 9648
rect 22100 9664 22152 9716
rect 25320 9707 25372 9716
rect 25320 9673 25329 9707
rect 25329 9673 25363 9707
rect 25363 9673 25372 9707
rect 25320 9664 25372 9673
rect 26148 9707 26200 9716
rect 26148 9673 26157 9707
rect 26157 9673 26191 9707
rect 26191 9673 26200 9707
rect 26148 9664 26200 9673
rect 29368 9664 29420 9716
rect 14096 9460 14148 9512
rect 16948 9528 17000 9580
rect 18696 9528 18748 9580
rect 19156 9571 19208 9580
rect 19156 9537 19165 9571
rect 19165 9537 19199 9571
rect 19199 9537 19208 9571
rect 19156 9528 19208 9537
rect 21548 9528 21600 9580
rect 21916 9571 21968 9580
rect 21916 9537 21925 9571
rect 21925 9537 21959 9571
rect 21959 9537 21968 9571
rect 22376 9596 22428 9648
rect 23204 9596 23256 9648
rect 25872 9596 25924 9648
rect 21916 9528 21968 9537
rect 22744 9528 22796 9580
rect 24952 9528 25004 9580
rect 23112 9460 23164 9512
rect 25412 9460 25464 9512
rect 8208 9324 8260 9376
rect 15660 9392 15712 9444
rect 16028 9392 16080 9444
rect 10140 9367 10192 9376
rect 10140 9333 10149 9367
rect 10149 9333 10183 9367
rect 10183 9333 10192 9367
rect 10140 9324 10192 9333
rect 11796 9367 11848 9376
rect 11796 9333 11805 9367
rect 11805 9333 11839 9367
rect 11839 9333 11848 9367
rect 11796 9324 11848 9333
rect 12992 9324 13044 9376
rect 13268 9367 13320 9376
rect 13268 9333 13277 9367
rect 13277 9333 13311 9367
rect 13311 9333 13320 9367
rect 13268 9324 13320 9333
rect 13360 9324 13412 9376
rect 19340 9324 19392 9376
rect 22560 9324 22612 9376
rect 22836 9324 22888 9376
rect 25228 9324 25280 9376
rect 26332 9528 26384 9580
rect 26976 9571 27028 9580
rect 26976 9537 26985 9571
rect 26985 9537 27019 9571
rect 27019 9537 27028 9571
rect 26976 9528 27028 9537
rect 28908 9596 28960 9648
rect 30380 9596 30432 9648
rect 32036 9596 32088 9648
rect 26608 9392 26660 9444
rect 31852 9528 31904 9580
rect 27528 9460 27580 9512
rect 29552 9460 29604 9512
rect 30288 9460 30340 9512
rect 31116 9503 31168 9512
rect 31116 9469 31125 9503
rect 31125 9469 31159 9503
rect 31159 9469 31168 9503
rect 31116 9460 31168 9469
rect 27252 9367 27304 9376
rect 27252 9333 27261 9367
rect 27261 9333 27295 9367
rect 27295 9333 27304 9367
rect 27252 9324 27304 9333
rect 32220 9367 32272 9376
rect 32220 9333 32229 9367
rect 32229 9333 32263 9367
rect 32263 9333 32272 9367
rect 32220 9324 32272 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 9128 9120 9180 9172
rect 8944 9052 8996 9104
rect 16028 9120 16080 9172
rect 16212 9163 16264 9172
rect 16212 9129 16221 9163
rect 16221 9129 16255 9163
rect 16255 9129 16264 9163
rect 16212 9120 16264 9129
rect 18696 9163 18748 9172
rect 18696 9129 18705 9163
rect 18705 9129 18739 9163
rect 18739 9129 18748 9163
rect 18696 9120 18748 9129
rect 21548 9163 21600 9172
rect 13912 9052 13964 9104
rect 21548 9129 21557 9163
rect 21557 9129 21591 9163
rect 21591 9129 21600 9163
rect 21548 9120 21600 9129
rect 22100 9120 22152 9172
rect 33140 9163 33192 9172
rect 33140 9129 33149 9163
rect 33149 9129 33183 9163
rect 33183 9129 33192 9163
rect 33140 9120 33192 9129
rect 7932 8984 7984 9036
rect 9588 8984 9640 9036
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 9128 8959 9180 8968
rect 9128 8925 9137 8959
rect 9137 8925 9171 8959
rect 9171 8925 9180 8959
rect 9128 8916 9180 8925
rect 11520 8984 11572 9036
rect 11796 8916 11848 8968
rect 12348 8916 12400 8968
rect 18328 9027 18380 9036
rect 18328 8993 18337 9027
rect 18337 8993 18371 9027
rect 18371 8993 18380 9027
rect 18328 8984 18380 8993
rect 14832 8959 14884 8968
rect 14832 8925 14841 8959
rect 14841 8925 14875 8959
rect 14875 8925 14884 8959
rect 14832 8916 14884 8925
rect 10140 8848 10192 8900
rect 13268 8848 13320 8900
rect 16948 8916 17000 8968
rect 18512 8959 18564 8968
rect 18512 8925 18521 8959
rect 18521 8925 18555 8959
rect 18555 8925 18564 8959
rect 18512 8916 18564 8925
rect 19248 8959 19300 8968
rect 19248 8925 19257 8959
rect 19257 8925 19291 8959
rect 19291 8925 19300 8959
rect 19248 8916 19300 8925
rect 19340 8916 19392 8968
rect 21364 8959 21416 8968
rect 16672 8848 16724 8900
rect 21364 8925 21373 8959
rect 21373 8925 21407 8959
rect 21407 8925 21416 8959
rect 21364 8916 21416 8925
rect 22836 8984 22888 9036
rect 25412 8984 25464 9036
rect 26884 8984 26936 9036
rect 21456 8848 21508 8900
rect 22192 8891 22244 8900
rect 22192 8857 22201 8891
rect 22201 8857 22235 8891
rect 22235 8857 22244 8891
rect 22192 8848 22244 8857
rect 22284 8891 22336 8900
rect 22284 8857 22293 8891
rect 22293 8857 22327 8891
rect 22327 8857 22336 8891
rect 22284 8848 22336 8857
rect 23020 8959 23072 8968
rect 23020 8925 23029 8959
rect 23029 8925 23063 8959
rect 23063 8925 23072 8959
rect 23020 8916 23072 8925
rect 23204 8916 23256 8968
rect 26240 8916 26292 8968
rect 29000 8916 29052 8968
rect 32588 8916 32640 8968
rect 25136 8848 25188 8900
rect 25320 8848 25372 8900
rect 27252 8848 27304 8900
rect 32220 8848 32272 8900
rect 34612 8848 34664 8900
rect 9680 8780 9732 8832
rect 9864 8780 9916 8832
rect 15476 8823 15528 8832
rect 15476 8789 15485 8823
rect 15485 8789 15519 8823
rect 15519 8789 15528 8823
rect 15476 8780 15528 8789
rect 18604 8780 18656 8832
rect 22468 8780 22520 8832
rect 22652 8780 22704 8832
rect 24768 8780 24820 8832
rect 24860 8780 24912 8832
rect 26516 8780 26568 8832
rect 27804 8780 27856 8832
rect 27988 8823 28040 8832
rect 27988 8789 27997 8823
rect 27997 8789 28031 8823
rect 28031 8789 28040 8823
rect 27988 8780 28040 8789
rect 30288 8780 30340 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 9128 8576 9180 8628
rect 4620 8508 4672 8560
rect 11520 8576 11572 8628
rect 13912 8576 13964 8628
rect 14096 8619 14148 8628
rect 14096 8585 14105 8619
rect 14105 8585 14139 8619
rect 14139 8585 14148 8619
rect 14096 8576 14148 8585
rect 16212 8576 16264 8628
rect 17960 8576 18012 8628
rect 18512 8576 18564 8628
rect 20536 8576 20588 8628
rect 24952 8619 25004 8628
rect 24952 8585 24961 8619
rect 24961 8585 24995 8619
rect 24995 8585 25004 8619
rect 24952 8576 25004 8585
rect 25596 8619 25648 8628
rect 25596 8585 25605 8619
rect 25605 8585 25639 8619
rect 25639 8585 25648 8619
rect 25596 8576 25648 8585
rect 8208 8483 8260 8492
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 8576 8483 8628 8492
rect 8576 8449 8585 8483
rect 8585 8449 8619 8483
rect 8619 8449 8628 8483
rect 8576 8440 8628 8449
rect 8760 8440 8812 8492
rect 9220 8483 9272 8492
rect 9220 8449 9229 8483
rect 9229 8449 9263 8483
rect 9263 8449 9272 8483
rect 9220 8440 9272 8449
rect 9864 8372 9916 8424
rect 11796 8483 11848 8492
rect 11796 8449 11805 8483
rect 11805 8449 11839 8483
rect 11839 8449 11848 8483
rect 13544 8508 13596 8560
rect 11796 8440 11848 8449
rect 12072 8372 12124 8424
rect 7472 8279 7524 8288
rect 7472 8245 7481 8279
rect 7481 8245 7515 8279
rect 7515 8245 7524 8279
rect 7472 8236 7524 8245
rect 8392 8304 8444 8356
rect 12992 8483 13044 8492
rect 12992 8449 13026 8483
rect 13026 8449 13044 8483
rect 12992 8440 13044 8449
rect 16120 8508 16172 8560
rect 15476 8440 15528 8492
rect 18788 8551 18840 8560
rect 18788 8517 18797 8551
rect 18797 8517 18831 8551
rect 18831 8517 18840 8551
rect 18788 8508 18840 8517
rect 23296 8508 23348 8560
rect 23480 8508 23532 8560
rect 24676 8551 24728 8560
rect 24676 8517 24685 8551
rect 24685 8517 24719 8551
rect 24719 8517 24728 8551
rect 24676 8508 24728 8517
rect 15844 8372 15896 8424
rect 17776 8483 17828 8492
rect 17776 8449 17785 8483
rect 17785 8449 17819 8483
rect 17819 8449 17828 8483
rect 17776 8440 17828 8449
rect 18604 8440 18656 8492
rect 18696 8483 18748 8492
rect 18696 8449 18705 8483
rect 18705 8449 18739 8483
rect 18739 8449 18748 8483
rect 18696 8440 18748 8449
rect 19616 8440 19668 8492
rect 21640 8440 21692 8492
rect 21732 8440 21784 8492
rect 22652 8440 22704 8492
rect 24216 8440 24268 8492
rect 24492 8440 24544 8492
rect 24768 8483 24820 8492
rect 24768 8449 24777 8483
rect 24777 8449 24811 8483
rect 24811 8449 24820 8483
rect 25412 8483 25464 8492
rect 24768 8440 24820 8449
rect 25412 8449 25421 8483
rect 25421 8449 25455 8483
rect 25455 8449 25464 8483
rect 25412 8440 25464 8449
rect 26424 8483 26476 8492
rect 26424 8449 26433 8483
rect 26433 8449 26467 8483
rect 26467 8449 26476 8483
rect 26424 8440 26476 8449
rect 27528 8508 27580 8560
rect 27712 8508 27764 8560
rect 20168 8415 20220 8424
rect 15936 8304 15988 8356
rect 20168 8381 20177 8415
rect 20177 8381 20211 8415
rect 20211 8381 20220 8415
rect 20168 8372 20220 8381
rect 21456 8372 21508 8424
rect 22284 8372 22336 8424
rect 27804 8440 27856 8492
rect 18696 8304 18748 8356
rect 21272 8304 21324 8356
rect 22376 8304 22428 8356
rect 9404 8236 9456 8288
rect 11796 8236 11848 8288
rect 12164 8236 12216 8288
rect 14924 8236 14976 8288
rect 15292 8236 15344 8288
rect 18512 8236 18564 8288
rect 21456 8236 21508 8288
rect 22284 8236 22336 8288
rect 23112 8236 23164 8288
rect 30104 8440 30156 8492
rect 32312 8440 32364 8492
rect 34612 8483 34664 8492
rect 34612 8449 34621 8483
rect 34621 8449 34655 8483
rect 34655 8449 34664 8483
rect 34612 8440 34664 8449
rect 34796 8483 34848 8492
rect 34796 8449 34805 8483
rect 34805 8449 34839 8483
rect 34839 8449 34848 8483
rect 34796 8440 34848 8449
rect 30288 8372 30340 8424
rect 32588 8415 32640 8424
rect 32588 8381 32597 8415
rect 32597 8381 32631 8415
rect 32631 8381 32640 8415
rect 32588 8372 32640 8381
rect 25044 8236 25096 8288
rect 26792 8236 26844 8288
rect 33968 8347 34020 8356
rect 33968 8313 33977 8347
rect 33977 8313 34011 8347
rect 34011 8313 34020 8347
rect 33968 8304 34020 8313
rect 29828 8279 29880 8288
rect 29828 8245 29837 8279
rect 29837 8245 29871 8279
rect 29871 8245 29880 8279
rect 29828 8236 29880 8245
rect 29920 8236 29972 8288
rect 33232 8236 33284 8288
rect 34520 8236 34572 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 8208 8075 8260 8084
rect 8208 8041 8217 8075
rect 8217 8041 8251 8075
rect 8251 8041 8260 8075
rect 8208 8032 8260 8041
rect 11060 8075 11112 8084
rect 11060 8041 11069 8075
rect 11069 8041 11103 8075
rect 11103 8041 11112 8075
rect 11060 8032 11112 8041
rect 11980 8075 12032 8084
rect 11980 8041 11989 8075
rect 11989 8041 12023 8075
rect 12023 8041 12032 8075
rect 11980 8032 12032 8041
rect 14832 8032 14884 8084
rect 15660 8032 15712 8084
rect 8576 7896 8628 7948
rect 12164 7964 12216 8016
rect 12992 7964 13044 8016
rect 15568 8007 15620 8016
rect 15568 7973 15577 8007
rect 15577 7973 15611 8007
rect 15611 7973 15620 8007
rect 15568 7964 15620 7973
rect 16672 8007 16724 8016
rect 16672 7973 16681 8007
rect 16681 7973 16715 8007
rect 16715 7973 16724 8007
rect 16672 7964 16724 7973
rect 19156 8032 19208 8084
rect 21364 8032 21416 8084
rect 22744 8032 22796 8084
rect 25136 8075 25188 8084
rect 25136 8041 25145 8075
rect 25145 8041 25179 8075
rect 25179 8041 25188 8075
rect 25136 8032 25188 8041
rect 28632 8032 28684 8084
rect 29184 8032 29236 8084
rect 7932 7828 7984 7880
rect 9680 7871 9732 7880
rect 9680 7837 9689 7871
rect 9689 7837 9723 7871
rect 9723 7837 9732 7871
rect 9680 7828 9732 7837
rect 9864 7871 9916 7880
rect 9864 7837 9873 7871
rect 9873 7837 9907 7871
rect 9907 7837 9916 7871
rect 9864 7828 9916 7837
rect 12348 7896 12400 7948
rect 11796 7871 11848 7880
rect 7472 7760 7524 7812
rect 11796 7837 11805 7871
rect 11805 7837 11839 7871
rect 11839 7837 11848 7871
rect 11796 7828 11848 7837
rect 15844 7896 15896 7948
rect 16212 7896 16264 7948
rect 17960 7896 18012 7948
rect 18328 7939 18380 7948
rect 18328 7905 18337 7939
rect 18337 7905 18371 7939
rect 18371 7905 18380 7939
rect 18328 7896 18380 7905
rect 18880 7896 18932 7948
rect 19156 7896 19208 7948
rect 19616 7896 19668 7948
rect 9496 7692 9548 7744
rect 14924 7828 14976 7880
rect 15476 7871 15528 7880
rect 14556 7760 14608 7812
rect 15476 7837 15485 7871
rect 15485 7837 15519 7871
rect 15519 7837 15528 7871
rect 15476 7828 15528 7837
rect 18512 7871 18564 7880
rect 18512 7837 18521 7871
rect 18521 7837 18555 7871
rect 18555 7837 18564 7871
rect 18512 7828 18564 7837
rect 20720 7828 20772 7880
rect 21732 7828 21784 7880
rect 23296 7896 23348 7948
rect 26240 7896 26292 7948
rect 22284 7871 22336 7880
rect 22284 7837 22293 7871
rect 22293 7837 22327 7871
rect 22327 7837 22336 7871
rect 22284 7828 22336 7837
rect 22468 7871 22520 7880
rect 22468 7837 22477 7871
rect 22477 7837 22511 7871
rect 22511 7837 22520 7871
rect 22468 7828 22520 7837
rect 23204 7871 23256 7880
rect 23204 7837 23213 7871
rect 23213 7837 23247 7871
rect 23247 7837 23256 7871
rect 23204 7828 23256 7837
rect 25228 7828 25280 7880
rect 15292 7692 15344 7744
rect 19432 7760 19484 7812
rect 18052 7692 18104 7744
rect 18512 7692 18564 7744
rect 23296 7760 23348 7812
rect 23480 7760 23532 7812
rect 26792 7896 26844 7948
rect 29920 7964 29972 8016
rect 26884 7871 26936 7880
rect 26884 7837 26893 7871
rect 26893 7837 26927 7871
rect 26927 7837 26936 7871
rect 26884 7828 26936 7837
rect 27528 7871 27580 7880
rect 27528 7837 27537 7871
rect 27537 7837 27571 7871
rect 27571 7837 27580 7871
rect 27528 7828 27580 7837
rect 28356 7828 28408 7880
rect 29644 7828 29696 7880
rect 33232 8032 33284 8084
rect 32312 8007 32364 8016
rect 32312 7973 32321 8007
rect 32321 7973 32355 8007
rect 32355 7973 32364 8007
rect 32312 7964 32364 7973
rect 32588 7964 32640 8016
rect 32680 7896 32732 7948
rect 27804 7803 27856 7812
rect 27804 7769 27838 7803
rect 27838 7769 27856 7803
rect 27804 7760 27856 7769
rect 28080 7760 28132 7812
rect 28908 7760 28960 7812
rect 29460 7760 29512 7812
rect 21272 7692 21324 7744
rect 23572 7692 23624 7744
rect 25320 7692 25372 7744
rect 27252 7692 27304 7744
rect 27712 7692 27764 7744
rect 33968 7828 34020 7880
rect 34520 7828 34572 7880
rect 37188 7828 37240 7880
rect 33140 7692 33192 7744
rect 34612 7692 34664 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 8392 7488 8444 7540
rect 9404 7531 9456 7540
rect 9404 7497 9413 7531
rect 9413 7497 9447 7531
rect 9447 7497 9456 7531
rect 9404 7488 9456 7497
rect 15476 7488 15528 7540
rect 8116 7352 8168 7404
rect 8300 7395 8352 7404
rect 8300 7361 8309 7395
rect 8309 7361 8343 7395
rect 8343 7361 8352 7395
rect 8300 7352 8352 7361
rect 8576 7420 8628 7472
rect 12992 7463 13044 7472
rect 12992 7429 13001 7463
rect 13001 7429 13035 7463
rect 13035 7429 13044 7463
rect 12992 7420 13044 7429
rect 12716 7395 12768 7404
rect 12716 7361 12725 7395
rect 12725 7361 12759 7395
rect 12759 7361 12768 7395
rect 12716 7352 12768 7361
rect 8944 7284 8996 7336
rect 11060 7284 11112 7336
rect 12072 7216 12124 7268
rect 13452 7352 13504 7404
rect 17224 7352 17276 7404
rect 18052 7352 18104 7404
rect 21272 7463 21324 7472
rect 21272 7429 21281 7463
rect 21281 7429 21315 7463
rect 21315 7429 21324 7463
rect 21272 7420 21324 7429
rect 21916 7420 21968 7472
rect 23480 7420 23532 7472
rect 24860 7420 24912 7472
rect 25412 7420 25464 7472
rect 26424 7420 26476 7472
rect 28356 7420 28408 7472
rect 30012 7420 30064 7472
rect 33140 7420 33192 7472
rect 34796 7488 34848 7540
rect 34336 7420 34388 7472
rect 20536 7395 20588 7404
rect 13544 7327 13596 7336
rect 13544 7293 13553 7327
rect 13553 7293 13587 7327
rect 13587 7293 13596 7327
rect 13544 7284 13596 7293
rect 17960 7284 18012 7336
rect 20536 7361 20545 7395
rect 20545 7361 20579 7395
rect 20579 7361 20588 7395
rect 20536 7352 20588 7361
rect 22468 7352 22520 7404
rect 23020 7352 23072 7404
rect 23940 7395 23992 7404
rect 23940 7361 23949 7395
rect 23949 7361 23983 7395
rect 23983 7361 23992 7395
rect 23940 7352 23992 7361
rect 26332 7395 26384 7404
rect 26332 7361 26341 7395
rect 26341 7361 26375 7395
rect 26375 7361 26384 7395
rect 26332 7352 26384 7361
rect 26884 7352 26936 7404
rect 22008 7284 22060 7336
rect 24952 7284 25004 7336
rect 25136 7327 25188 7336
rect 25136 7293 25145 7327
rect 25145 7293 25179 7327
rect 25179 7293 25188 7327
rect 25136 7284 25188 7293
rect 26976 7327 27028 7336
rect 26976 7293 26985 7327
rect 26985 7293 27019 7327
rect 27019 7293 27028 7327
rect 26976 7284 27028 7293
rect 27252 7352 27304 7404
rect 27988 7395 28040 7404
rect 27988 7361 27997 7395
rect 27997 7361 28031 7395
rect 28031 7361 28040 7395
rect 27988 7352 28040 7361
rect 28540 7352 28592 7404
rect 29828 7352 29880 7404
rect 30380 7395 30432 7404
rect 30380 7361 30414 7395
rect 30414 7361 30432 7395
rect 30380 7352 30432 7361
rect 34612 7395 34664 7404
rect 34612 7361 34621 7395
rect 34621 7361 34655 7395
rect 34655 7361 34664 7395
rect 34612 7352 34664 7361
rect 37924 7420 37976 7472
rect 13360 7148 13412 7200
rect 16672 7148 16724 7200
rect 19432 7216 19484 7268
rect 19524 7148 19576 7200
rect 20352 7191 20404 7200
rect 20352 7157 20361 7191
rect 20361 7157 20395 7191
rect 20395 7157 20404 7191
rect 20352 7148 20404 7157
rect 23020 7148 23072 7200
rect 25320 7148 25372 7200
rect 27804 7191 27856 7200
rect 27804 7157 27813 7191
rect 27813 7157 27847 7191
rect 27847 7157 27856 7191
rect 27804 7148 27856 7157
rect 28356 7148 28408 7200
rect 28724 7148 28776 7200
rect 29000 7191 29052 7200
rect 29000 7157 29009 7191
rect 29009 7157 29043 7191
rect 29043 7157 29052 7191
rect 29000 7148 29052 7157
rect 29460 7191 29512 7200
rect 29460 7157 29469 7191
rect 29469 7157 29503 7191
rect 29503 7157 29512 7191
rect 29460 7148 29512 7157
rect 29644 7216 29696 7268
rect 33140 7284 33192 7336
rect 35440 7216 35492 7268
rect 31484 7191 31536 7200
rect 31484 7157 31493 7191
rect 31493 7157 31527 7191
rect 31527 7157 31536 7191
rect 31484 7148 31536 7157
rect 32680 7191 32732 7200
rect 32680 7157 32689 7191
rect 32689 7157 32723 7191
rect 32723 7157 32732 7191
rect 32680 7148 32732 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 18052 6987 18104 6996
rect 18052 6953 18061 6987
rect 18061 6953 18095 6987
rect 18095 6953 18104 6987
rect 18052 6944 18104 6953
rect 19432 6944 19484 6996
rect 9588 6808 9640 6860
rect 8944 6740 8996 6792
rect 8392 6672 8444 6724
rect 9312 6672 9364 6724
rect 9956 6672 10008 6724
rect 10600 6740 10652 6792
rect 12992 6808 13044 6860
rect 13452 6851 13504 6860
rect 13452 6817 13461 6851
rect 13461 6817 13495 6851
rect 13495 6817 13504 6851
rect 13452 6808 13504 6817
rect 16120 6851 16172 6860
rect 11980 6740 12032 6792
rect 13360 6783 13412 6792
rect 13360 6749 13369 6783
rect 13369 6749 13403 6783
rect 13403 6749 13412 6783
rect 13360 6740 13412 6749
rect 15476 6783 15528 6792
rect 11152 6672 11204 6724
rect 10416 6604 10468 6656
rect 12532 6647 12584 6656
rect 12532 6613 12541 6647
rect 12541 6613 12575 6647
rect 12575 6613 12584 6647
rect 12532 6604 12584 6613
rect 12900 6672 12952 6724
rect 15476 6749 15485 6783
rect 15485 6749 15519 6783
rect 15519 6749 15528 6783
rect 15476 6740 15528 6749
rect 16120 6817 16129 6851
rect 16129 6817 16163 6851
rect 16163 6817 16172 6851
rect 16120 6808 16172 6817
rect 18144 6808 18196 6860
rect 21364 6944 21416 6996
rect 22008 6944 22060 6996
rect 25136 6944 25188 6996
rect 26424 6944 26476 6996
rect 26976 6944 27028 6996
rect 27528 6944 27580 6996
rect 29000 6944 29052 6996
rect 31484 6944 31536 6996
rect 33968 6944 34020 6996
rect 24676 6876 24728 6928
rect 28080 6876 28132 6928
rect 22376 6851 22428 6860
rect 22376 6817 22385 6851
rect 22385 6817 22419 6851
rect 22419 6817 22428 6851
rect 22376 6808 22428 6817
rect 24124 6808 24176 6860
rect 17960 6740 18012 6792
rect 18236 6783 18288 6792
rect 18236 6749 18245 6783
rect 18245 6749 18279 6783
rect 18279 6749 18288 6783
rect 18236 6740 18288 6749
rect 19524 6783 19576 6792
rect 19524 6749 19533 6783
rect 19533 6749 19567 6783
rect 19567 6749 19576 6783
rect 19524 6740 19576 6749
rect 22100 6740 22152 6792
rect 22284 6740 22336 6792
rect 24676 6740 24728 6792
rect 26240 6740 26292 6792
rect 32312 6808 32364 6860
rect 35808 6808 35860 6860
rect 14280 6604 14332 6656
rect 16856 6604 16908 6656
rect 20352 6672 20404 6724
rect 22836 6672 22888 6724
rect 23296 6672 23348 6724
rect 20628 6604 20680 6656
rect 21824 6604 21876 6656
rect 22192 6604 22244 6656
rect 24492 6672 24544 6724
rect 25044 6647 25096 6656
rect 25044 6613 25053 6647
rect 25053 6613 25087 6647
rect 25087 6613 25096 6647
rect 25044 6604 25096 6613
rect 26056 6672 26108 6724
rect 29184 6740 29236 6792
rect 29920 6783 29972 6792
rect 29920 6749 29929 6783
rect 29929 6749 29963 6783
rect 29963 6749 29972 6783
rect 29920 6740 29972 6749
rect 30288 6740 30340 6792
rect 30748 6783 30800 6792
rect 30748 6749 30757 6783
rect 30757 6749 30791 6783
rect 30791 6749 30800 6783
rect 30748 6740 30800 6749
rect 31760 6783 31812 6792
rect 31760 6749 31769 6783
rect 31769 6749 31803 6783
rect 31803 6749 31812 6783
rect 31760 6740 31812 6749
rect 32128 6740 32180 6792
rect 32680 6783 32732 6792
rect 32680 6749 32714 6783
rect 32714 6749 32732 6783
rect 32680 6740 32732 6749
rect 34612 6740 34664 6792
rect 27620 6672 27672 6724
rect 28724 6672 28776 6724
rect 29276 6672 29328 6724
rect 30104 6647 30156 6656
rect 30104 6613 30113 6647
rect 30113 6613 30147 6647
rect 30147 6613 30156 6647
rect 30104 6604 30156 6613
rect 30472 6604 30524 6656
rect 33324 6604 33376 6656
rect 34796 6604 34848 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 7748 6307 7800 6316
rect 7748 6273 7757 6307
rect 7757 6273 7791 6307
rect 7791 6273 7800 6307
rect 7748 6264 7800 6273
rect 8392 6400 8444 6452
rect 9128 6400 9180 6452
rect 8484 6332 8536 6384
rect 9588 6332 9640 6384
rect 10692 6375 10744 6384
rect 10692 6341 10701 6375
rect 10701 6341 10735 6375
rect 10735 6341 10744 6375
rect 10692 6332 10744 6341
rect 12532 6332 12584 6384
rect 13176 6400 13228 6452
rect 14556 6400 14608 6452
rect 15108 6443 15160 6452
rect 15108 6409 15117 6443
rect 15117 6409 15151 6443
rect 15151 6409 15160 6443
rect 15108 6400 15160 6409
rect 13820 6332 13872 6384
rect 10416 6307 10468 6316
rect 10416 6273 10425 6307
rect 10425 6273 10459 6307
rect 10459 6273 10468 6307
rect 10416 6264 10468 6273
rect 11796 6264 11848 6316
rect 12900 6264 12952 6316
rect 11612 6196 11664 6248
rect 10784 6060 10836 6112
rect 12808 6196 12860 6248
rect 15476 6332 15528 6384
rect 17592 6400 17644 6452
rect 18604 6400 18656 6452
rect 18696 6400 18748 6452
rect 20168 6400 20220 6452
rect 20536 6400 20588 6452
rect 20628 6400 20680 6452
rect 18144 6332 18196 6384
rect 14096 6264 14148 6316
rect 15016 6264 15068 6316
rect 14740 6196 14792 6248
rect 16672 6239 16724 6248
rect 16672 6205 16681 6239
rect 16681 6205 16715 6239
rect 16715 6205 16724 6239
rect 16672 6196 16724 6205
rect 16856 6239 16908 6248
rect 16856 6205 16865 6239
rect 16865 6205 16899 6239
rect 16899 6205 16908 6239
rect 16856 6196 16908 6205
rect 17132 6264 17184 6316
rect 17408 6264 17460 6316
rect 18236 6264 18288 6316
rect 18696 6307 18748 6316
rect 18696 6273 18705 6307
rect 18705 6273 18739 6307
rect 18739 6273 18748 6307
rect 18696 6264 18748 6273
rect 21364 6332 21416 6384
rect 22468 6400 22520 6452
rect 22836 6443 22888 6452
rect 22836 6409 22845 6443
rect 22845 6409 22879 6443
rect 22879 6409 22888 6443
rect 22836 6400 22888 6409
rect 26240 6400 26292 6452
rect 27068 6400 27120 6452
rect 28080 6443 28132 6452
rect 28080 6409 28089 6443
rect 28089 6409 28123 6443
rect 28123 6409 28132 6443
rect 28080 6400 28132 6409
rect 21088 6307 21140 6316
rect 17316 6196 17368 6248
rect 18604 6196 18656 6248
rect 14188 6128 14240 6180
rect 16948 6171 17000 6180
rect 16948 6137 16957 6171
rect 16957 6137 16991 6171
rect 16991 6137 17000 6171
rect 16948 6128 17000 6137
rect 18880 6128 18932 6180
rect 12440 6060 12492 6112
rect 12716 6060 12768 6112
rect 13912 6060 13964 6112
rect 14648 6060 14700 6112
rect 18696 6060 18748 6112
rect 21088 6273 21097 6307
rect 21097 6273 21131 6307
rect 21131 6273 21140 6307
rect 21088 6264 21140 6273
rect 21824 6307 21876 6316
rect 21824 6273 21833 6307
rect 21833 6273 21867 6307
rect 21867 6273 21876 6307
rect 21824 6264 21876 6273
rect 22928 6332 22980 6384
rect 24860 6332 24912 6384
rect 26976 6332 27028 6384
rect 30380 6400 30432 6452
rect 31024 6400 31076 6452
rect 23020 6307 23072 6316
rect 21732 6060 21784 6112
rect 23020 6273 23029 6307
rect 23029 6273 23063 6307
rect 23063 6273 23072 6307
rect 23020 6264 23072 6273
rect 23756 6307 23808 6316
rect 23756 6273 23765 6307
rect 23765 6273 23799 6307
rect 23799 6273 23808 6307
rect 23756 6264 23808 6273
rect 25044 6307 25096 6316
rect 25044 6273 25053 6307
rect 25053 6273 25087 6307
rect 25087 6273 25096 6307
rect 25044 6264 25096 6273
rect 25320 6307 25372 6316
rect 25320 6273 25354 6307
rect 25354 6273 25372 6307
rect 25320 6264 25372 6273
rect 27068 6307 27120 6316
rect 27068 6273 27077 6307
rect 27077 6273 27111 6307
rect 27111 6273 27120 6307
rect 27068 6264 27120 6273
rect 22468 6196 22520 6248
rect 22744 6196 22796 6248
rect 24676 6196 24728 6248
rect 27436 6307 27488 6316
rect 27436 6273 27445 6307
rect 27445 6273 27479 6307
rect 27479 6273 27488 6307
rect 27436 6264 27488 6273
rect 27620 6264 27672 6316
rect 29000 6264 29052 6316
rect 29276 6264 29328 6316
rect 29460 6307 29512 6316
rect 29460 6273 29469 6307
rect 29469 6273 29503 6307
rect 29503 6273 29512 6307
rect 29460 6264 29512 6273
rect 30748 6332 30800 6384
rect 31208 6332 31260 6384
rect 32772 6400 32824 6452
rect 29920 6264 29972 6316
rect 30472 6307 30524 6316
rect 30472 6273 30481 6307
rect 30481 6273 30515 6307
rect 30515 6273 30524 6307
rect 30472 6264 30524 6273
rect 31116 6307 31168 6316
rect 31116 6273 31125 6307
rect 31125 6273 31159 6307
rect 31159 6273 31168 6307
rect 31116 6264 31168 6273
rect 32956 6264 33008 6316
rect 33324 6264 33376 6316
rect 34060 6307 34112 6316
rect 23848 6060 23900 6112
rect 31944 6196 31996 6248
rect 32404 6239 32456 6248
rect 32404 6205 32413 6239
rect 32413 6205 32447 6239
rect 32447 6205 32456 6239
rect 32404 6196 32456 6205
rect 34060 6273 34069 6307
rect 34069 6273 34103 6307
rect 34103 6273 34112 6307
rect 34060 6264 34112 6273
rect 35624 6196 35676 6248
rect 31668 6128 31720 6180
rect 26516 6060 26568 6112
rect 28724 6060 28776 6112
rect 31300 6060 31352 6112
rect 33416 6128 33468 6180
rect 33140 6060 33192 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 7748 5856 7800 5908
rect 9956 5899 10008 5908
rect 9956 5865 9965 5899
rect 9965 5865 9999 5899
rect 9999 5865 10008 5899
rect 9956 5856 10008 5865
rect 9588 5788 9640 5840
rect 16948 5856 17000 5908
rect 17776 5899 17828 5908
rect 17776 5865 17785 5899
rect 17785 5865 17819 5899
rect 17819 5865 17828 5899
rect 17776 5856 17828 5865
rect 9128 5763 9180 5772
rect 9128 5729 9137 5763
rect 9137 5729 9171 5763
rect 9171 5729 9180 5763
rect 9128 5720 9180 5729
rect 5540 5652 5592 5704
rect 10600 5695 10652 5704
rect 10600 5661 10609 5695
rect 10609 5661 10643 5695
rect 10643 5661 10652 5695
rect 10600 5652 10652 5661
rect 10784 5695 10836 5704
rect 10784 5661 10793 5695
rect 10793 5661 10827 5695
rect 10827 5661 10836 5695
rect 10784 5652 10836 5661
rect 12716 5788 12768 5840
rect 14648 5788 14700 5840
rect 15752 5788 15804 5840
rect 12992 5763 13044 5772
rect 12992 5729 13001 5763
rect 13001 5729 13035 5763
rect 13035 5729 13044 5763
rect 12992 5720 13044 5729
rect 16120 5720 16172 5772
rect 11612 5695 11664 5704
rect 11612 5661 11621 5695
rect 11621 5661 11655 5695
rect 11655 5661 11664 5695
rect 11612 5652 11664 5661
rect 11888 5652 11940 5704
rect 10416 5584 10468 5636
rect 12808 5652 12860 5704
rect 14648 5695 14700 5704
rect 14648 5661 14657 5695
rect 14657 5661 14691 5695
rect 14691 5661 14700 5695
rect 14648 5652 14700 5661
rect 11428 5516 11480 5568
rect 16212 5584 16264 5636
rect 16764 5652 16816 5704
rect 17316 5695 17368 5704
rect 17316 5661 17325 5695
rect 17325 5661 17359 5695
rect 17359 5661 17368 5695
rect 17316 5652 17368 5661
rect 19432 5856 19484 5908
rect 20168 5856 20220 5908
rect 21732 5899 21784 5908
rect 21732 5865 21741 5899
rect 21741 5865 21775 5899
rect 21775 5865 21784 5899
rect 21732 5856 21784 5865
rect 26332 5856 26384 5908
rect 21088 5788 21140 5840
rect 24768 5788 24820 5840
rect 25136 5788 25188 5840
rect 27620 5856 27672 5908
rect 27896 5856 27948 5908
rect 28724 5856 28776 5908
rect 26884 5788 26936 5840
rect 19248 5763 19300 5772
rect 19248 5729 19257 5763
rect 19257 5729 19291 5763
rect 19291 5729 19300 5763
rect 19248 5720 19300 5729
rect 18880 5652 18932 5704
rect 23572 5720 23624 5772
rect 22560 5652 22612 5704
rect 24860 5720 24912 5772
rect 27436 5720 27488 5772
rect 28816 5788 28868 5840
rect 30012 5856 30064 5908
rect 34704 5856 34756 5908
rect 35808 5856 35860 5908
rect 37924 5899 37976 5908
rect 37924 5865 37933 5899
rect 37933 5865 37967 5899
rect 37967 5865 37976 5899
rect 37924 5856 37976 5865
rect 24400 5695 24452 5704
rect 24400 5661 24409 5695
rect 24409 5661 24443 5695
rect 24443 5661 24452 5695
rect 24400 5652 24452 5661
rect 18604 5584 18656 5636
rect 19340 5584 19392 5636
rect 20536 5584 20588 5636
rect 11980 5559 12032 5568
rect 11980 5525 11989 5559
rect 11989 5525 12023 5559
rect 12023 5525 12032 5559
rect 11980 5516 12032 5525
rect 15476 5516 15528 5568
rect 16488 5559 16540 5568
rect 16488 5525 16497 5559
rect 16497 5525 16531 5559
rect 16531 5525 16540 5559
rect 16488 5516 16540 5525
rect 18972 5516 19024 5568
rect 19984 5516 20036 5568
rect 20352 5516 20404 5568
rect 21824 5584 21876 5636
rect 23940 5584 23992 5636
rect 24768 5652 24820 5704
rect 26332 5695 26384 5704
rect 26332 5661 26341 5695
rect 26341 5661 26375 5695
rect 26375 5661 26384 5695
rect 26332 5652 26384 5661
rect 26516 5695 26568 5704
rect 26516 5661 26525 5695
rect 26525 5661 26559 5695
rect 26559 5661 26568 5695
rect 26516 5652 26568 5661
rect 26884 5652 26936 5704
rect 27712 5652 27764 5704
rect 30564 5788 30616 5840
rect 22284 5516 22336 5568
rect 26424 5584 26476 5636
rect 24492 5559 24544 5568
rect 24492 5525 24501 5559
rect 24501 5525 24535 5559
rect 24535 5525 24544 5559
rect 24492 5516 24544 5525
rect 26240 5516 26292 5568
rect 26792 5516 26844 5568
rect 29092 5584 29144 5636
rect 29920 5652 29972 5704
rect 32312 5695 32364 5704
rect 29552 5516 29604 5568
rect 29736 5516 29788 5568
rect 30932 5584 30984 5636
rect 32312 5661 32321 5695
rect 32321 5661 32355 5695
rect 32355 5661 32364 5695
rect 32312 5652 32364 5661
rect 30380 5516 30432 5568
rect 31116 5516 31168 5568
rect 32128 5516 32180 5568
rect 39028 5652 39080 5704
rect 34520 5584 34572 5636
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 9496 5355 9548 5364
rect 9496 5321 9505 5355
rect 9505 5321 9539 5355
rect 9539 5321 9548 5355
rect 9496 5312 9548 5321
rect 10508 5312 10560 5364
rect 11704 5355 11756 5364
rect 11704 5321 11713 5355
rect 11713 5321 11747 5355
rect 11747 5321 11756 5355
rect 11704 5312 11756 5321
rect 18788 5312 18840 5364
rect 20076 5312 20128 5364
rect 22192 5312 22244 5364
rect 8760 5244 8812 5296
rect 20168 5244 20220 5296
rect 10232 5176 10284 5228
rect 10508 5176 10560 5228
rect 11612 5176 11664 5228
rect 14004 5176 14056 5228
rect 17224 5219 17276 5228
rect 17224 5185 17233 5219
rect 17233 5185 17267 5219
rect 17267 5185 17276 5219
rect 17224 5176 17276 5185
rect 12440 5108 12492 5160
rect 13544 5108 13596 5160
rect 14648 5108 14700 5160
rect 16856 5108 16908 5160
rect 16304 5040 16356 5092
rect 17960 5176 18012 5228
rect 18420 5176 18472 5228
rect 19248 5176 19300 5228
rect 22560 5244 22612 5296
rect 19984 5108 20036 5160
rect 17776 5040 17828 5092
rect 19708 5040 19760 5092
rect 21272 5176 21324 5228
rect 23204 5176 23256 5228
rect 25044 5244 25096 5296
rect 24492 5176 24544 5228
rect 26240 5219 26292 5228
rect 26240 5185 26249 5219
rect 26249 5185 26283 5219
rect 26283 5185 26292 5219
rect 26240 5176 26292 5185
rect 26424 5219 26476 5228
rect 26424 5185 26433 5219
rect 26433 5185 26467 5219
rect 26467 5185 26476 5219
rect 26424 5176 26476 5185
rect 27528 5176 27580 5228
rect 29644 5244 29696 5296
rect 26976 5151 27028 5160
rect 20996 5040 21048 5092
rect 13544 4972 13596 5024
rect 14280 4972 14332 5024
rect 17316 5015 17368 5024
rect 17316 4981 17325 5015
rect 17325 4981 17359 5015
rect 17359 4981 17368 5015
rect 17316 4972 17368 4981
rect 18052 5015 18104 5024
rect 18052 4981 18061 5015
rect 18061 4981 18095 5015
rect 18095 4981 18104 5015
rect 18052 4972 18104 4981
rect 18972 4972 19024 5024
rect 20904 4972 20956 5024
rect 22008 4972 22060 5024
rect 23204 4972 23256 5024
rect 26976 5117 26985 5151
rect 26985 5117 27019 5151
rect 27019 5117 27028 5151
rect 26976 5108 27028 5117
rect 27988 5108 28040 5160
rect 30472 5176 30524 5228
rect 31944 5244 31996 5296
rect 34520 5312 34572 5364
rect 31852 5176 31904 5228
rect 34612 5219 34664 5228
rect 32128 5151 32180 5160
rect 32128 5117 32137 5151
rect 32137 5117 32171 5151
rect 32171 5117 32180 5151
rect 32128 5108 32180 5117
rect 31576 5040 31628 5092
rect 34612 5185 34621 5219
rect 34621 5185 34655 5219
rect 34655 5185 34664 5219
rect 34612 5176 34664 5185
rect 35348 5176 35400 5228
rect 37832 5219 37884 5228
rect 37832 5185 37841 5219
rect 37841 5185 37875 5219
rect 37875 5185 37884 5219
rect 37832 5176 37884 5185
rect 24584 4972 24636 5024
rect 25412 5015 25464 5024
rect 25412 4981 25421 5015
rect 25421 4981 25455 5015
rect 25455 4981 25464 5015
rect 25412 4972 25464 4981
rect 27620 4972 27672 5024
rect 28356 5015 28408 5024
rect 28356 4981 28365 5015
rect 28365 4981 28399 5015
rect 28399 4981 28408 5015
rect 28356 4972 28408 4981
rect 28816 4972 28868 5024
rect 30748 5015 30800 5024
rect 30748 4981 30757 5015
rect 30757 4981 30791 5015
rect 30791 4981 30800 5015
rect 30748 4972 30800 4981
rect 32404 4972 32456 5024
rect 39764 4972 39816 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 10416 4768 10468 4820
rect 11796 4700 11848 4752
rect 13912 4768 13964 4820
rect 17592 4768 17644 4820
rect 18972 4768 19024 4820
rect 19340 4811 19392 4820
rect 19340 4777 19349 4811
rect 19349 4777 19383 4811
rect 19383 4777 19392 4811
rect 19340 4768 19392 4777
rect 22008 4811 22060 4820
rect 22008 4777 22017 4811
rect 22017 4777 22051 4811
rect 22051 4777 22060 4811
rect 22008 4768 22060 4777
rect 24400 4768 24452 4820
rect 25412 4768 25464 4820
rect 26240 4768 26292 4820
rect 27620 4768 27672 4820
rect 27988 4811 28040 4820
rect 14188 4700 14240 4752
rect 14280 4675 14332 4684
rect 14280 4641 14289 4675
rect 14289 4641 14323 4675
rect 14323 4641 14332 4675
rect 14280 4632 14332 4641
rect 15476 4675 15528 4684
rect 15476 4641 15485 4675
rect 15485 4641 15519 4675
rect 15519 4641 15528 4675
rect 15476 4632 15528 4641
rect 9128 4564 9180 4616
rect 9312 4564 9364 4616
rect 10140 4564 10192 4616
rect 11244 4564 11296 4616
rect 12440 4564 12492 4616
rect 12624 4564 12676 4616
rect 14188 4564 14240 4616
rect 10600 4496 10652 4548
rect 15292 4539 15344 4548
rect 15292 4505 15301 4539
rect 15301 4505 15335 4539
rect 15335 4505 15344 4539
rect 15292 4496 15344 4505
rect 9128 4471 9180 4480
rect 9128 4437 9137 4471
rect 9137 4437 9171 4471
rect 9171 4437 9180 4471
rect 9128 4428 9180 4437
rect 11336 4471 11388 4480
rect 11336 4437 11345 4471
rect 11345 4437 11379 4471
rect 11379 4437 11388 4471
rect 11336 4428 11388 4437
rect 12072 4471 12124 4480
rect 12072 4437 12081 4471
rect 12081 4437 12115 4471
rect 12115 4437 12124 4471
rect 12072 4428 12124 4437
rect 12808 4428 12860 4480
rect 13360 4471 13412 4480
rect 13360 4437 13369 4471
rect 13369 4437 13403 4471
rect 13403 4437 13412 4471
rect 13360 4428 13412 4437
rect 20812 4700 20864 4752
rect 16212 4675 16264 4684
rect 16212 4641 16221 4675
rect 16221 4641 16255 4675
rect 16255 4641 16264 4675
rect 16212 4632 16264 4641
rect 16304 4607 16356 4616
rect 16304 4573 16313 4607
rect 16313 4573 16347 4607
rect 16347 4573 16356 4607
rect 16856 4607 16908 4616
rect 16304 4564 16356 4573
rect 16488 4496 16540 4548
rect 16856 4573 16865 4607
rect 16865 4573 16899 4607
rect 16899 4573 16908 4607
rect 16856 4564 16908 4573
rect 17868 4564 17920 4616
rect 19248 4607 19300 4616
rect 19248 4573 19257 4607
rect 19257 4573 19291 4607
rect 19291 4573 19300 4607
rect 19248 4564 19300 4573
rect 20904 4632 20956 4684
rect 21732 4675 21784 4684
rect 20076 4607 20128 4616
rect 16948 4428 17000 4480
rect 17316 4496 17368 4548
rect 20076 4573 20085 4607
rect 20085 4573 20119 4607
rect 20119 4573 20128 4607
rect 20076 4564 20128 4573
rect 21732 4641 21741 4675
rect 21741 4641 21775 4675
rect 21775 4641 21784 4675
rect 21732 4632 21784 4641
rect 22192 4632 22244 4684
rect 22008 4564 22060 4616
rect 22468 4564 22520 4616
rect 23940 4632 23992 4684
rect 24584 4675 24636 4684
rect 24584 4641 24593 4675
rect 24593 4641 24627 4675
rect 24627 4641 24636 4675
rect 24584 4632 24636 4641
rect 23664 4564 23716 4616
rect 27988 4777 27997 4811
rect 27997 4777 28031 4811
rect 28031 4777 28040 4811
rect 27988 4768 28040 4777
rect 28816 4811 28868 4820
rect 28816 4777 28825 4811
rect 28825 4777 28859 4811
rect 28859 4777 28868 4811
rect 28816 4768 28868 4777
rect 28908 4768 28960 4820
rect 32220 4768 32272 4820
rect 32404 4811 32456 4820
rect 32404 4777 32413 4811
rect 32413 4777 32447 4811
rect 32447 4777 32456 4811
rect 32404 4768 32456 4777
rect 33140 4768 33192 4820
rect 35716 4811 35768 4820
rect 35716 4777 35725 4811
rect 35725 4777 35759 4811
rect 35759 4777 35768 4811
rect 35716 4768 35768 4777
rect 37188 4811 37240 4820
rect 37188 4777 37197 4811
rect 37197 4777 37231 4811
rect 37231 4777 37240 4811
rect 37188 4768 37240 4777
rect 28724 4700 28776 4752
rect 31116 4700 31168 4752
rect 26332 4632 26384 4684
rect 25596 4607 25648 4616
rect 25596 4573 25605 4607
rect 25605 4573 25639 4607
rect 25639 4573 25648 4607
rect 25596 4564 25648 4573
rect 27528 4632 27580 4684
rect 26792 4607 26844 4616
rect 26792 4573 26801 4607
rect 26801 4573 26835 4607
rect 26835 4573 26844 4607
rect 26792 4564 26844 4573
rect 27436 4607 27488 4616
rect 27436 4573 27445 4607
rect 27445 4573 27479 4607
rect 27479 4573 27488 4607
rect 27896 4607 27948 4616
rect 27436 4564 27488 4573
rect 27896 4573 27905 4607
rect 27905 4573 27939 4607
rect 27939 4573 27948 4607
rect 27896 4564 27948 4573
rect 28724 4607 28776 4616
rect 28724 4573 28733 4607
rect 28733 4573 28767 4607
rect 28767 4573 28776 4607
rect 28724 4564 28776 4573
rect 28356 4496 28408 4548
rect 29644 4564 29696 4616
rect 31576 4564 31628 4616
rect 18236 4471 18288 4480
rect 18236 4437 18245 4471
rect 18245 4437 18279 4471
rect 18279 4437 18288 4471
rect 18236 4428 18288 4437
rect 19984 4428 20036 4480
rect 22192 4428 22244 4480
rect 22284 4428 22336 4480
rect 23480 4471 23532 4480
rect 23480 4437 23489 4471
rect 23489 4437 23523 4471
rect 23523 4437 23532 4471
rect 23480 4428 23532 4437
rect 25320 4428 25372 4480
rect 29460 4428 29512 4480
rect 30748 4496 30800 4548
rect 30564 4428 30616 4480
rect 30840 4428 30892 4480
rect 31852 4428 31904 4480
rect 32588 4632 32640 4684
rect 33508 4564 33560 4616
rect 34336 4564 34388 4616
rect 34704 4607 34756 4616
rect 34428 4496 34480 4548
rect 34704 4573 34713 4607
rect 34713 4573 34747 4607
rect 34747 4573 34756 4607
rect 34704 4564 34756 4573
rect 35072 4607 35124 4616
rect 35072 4573 35081 4607
rect 35081 4573 35115 4607
rect 35115 4573 35124 4607
rect 35072 4564 35124 4573
rect 35256 4564 35308 4616
rect 36544 4496 36596 4548
rect 37924 4496 37976 4548
rect 34520 4428 34572 4480
rect 38660 4428 38712 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 15200 4224 15252 4276
rect 15292 4224 15344 4276
rect 9128 4156 9180 4208
rect 11520 4199 11572 4208
rect 11520 4165 11529 4199
rect 11529 4165 11563 4199
rect 11563 4165 11572 4199
rect 11520 4156 11572 4165
rect 12808 4199 12860 4208
rect 12808 4165 12817 4199
rect 12817 4165 12851 4199
rect 12851 4165 12860 4199
rect 12808 4156 12860 4165
rect 14280 4156 14332 4208
rect 8484 4088 8536 4140
rect 9588 4088 9640 4140
rect 11336 4088 11388 4140
rect 12532 4131 12584 4140
rect 12532 4097 12541 4131
rect 12541 4097 12575 4131
rect 12575 4097 12584 4131
rect 12532 4088 12584 4097
rect 13912 4131 13964 4140
rect 10416 3995 10468 4004
rect 10416 3961 10425 3995
rect 10425 3961 10459 3995
rect 10459 3961 10468 3995
rect 10416 3952 10468 3961
rect 11152 4020 11204 4072
rect 11704 4020 11756 4072
rect 13912 4097 13921 4131
rect 13921 4097 13955 4131
rect 13955 4097 13964 4131
rect 13912 4088 13964 4097
rect 14648 4131 14700 4140
rect 1676 3884 1728 3936
rect 3056 3884 3108 3936
rect 8852 3884 8904 3936
rect 8944 3884 8996 3936
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 12716 3884 12768 3936
rect 13820 4020 13872 4072
rect 14004 4063 14056 4072
rect 14004 4029 14013 4063
rect 14013 4029 14047 4063
rect 14047 4029 14056 4063
rect 14004 4020 14056 4029
rect 14648 4097 14657 4131
rect 14657 4097 14691 4131
rect 14691 4097 14700 4131
rect 14648 4088 14700 4097
rect 16304 4156 16356 4208
rect 15660 4131 15712 4140
rect 15660 4097 15669 4131
rect 15669 4097 15703 4131
rect 15703 4097 15712 4131
rect 15660 4088 15712 4097
rect 17040 4088 17092 4140
rect 17776 4224 17828 4276
rect 19156 4224 19208 4276
rect 18236 4156 18288 4208
rect 21088 4224 21140 4276
rect 22008 4224 22060 4276
rect 24400 4224 24452 4276
rect 29552 4224 29604 4276
rect 18052 4088 18104 4140
rect 14924 4020 14976 4072
rect 13636 3952 13688 4004
rect 16764 4020 16816 4072
rect 18236 4020 18288 4072
rect 16396 3952 16448 4004
rect 17592 3995 17644 4004
rect 17592 3961 17601 3995
rect 17601 3961 17635 3995
rect 17635 3961 17644 3995
rect 17592 3952 17644 3961
rect 17776 3952 17828 4004
rect 18512 4088 18564 4140
rect 19248 4131 19300 4140
rect 19248 4097 19257 4131
rect 19257 4097 19291 4131
rect 19291 4097 19300 4131
rect 19248 4088 19300 4097
rect 22192 4156 22244 4208
rect 24768 4156 24820 4208
rect 26240 4156 26292 4208
rect 21088 4131 21140 4140
rect 19156 4063 19208 4072
rect 19156 4029 19165 4063
rect 19165 4029 19199 4063
rect 19199 4029 19208 4063
rect 19156 4020 19208 4029
rect 14464 3884 14516 3936
rect 15292 3884 15344 3936
rect 15476 3927 15528 3936
rect 15476 3893 15485 3927
rect 15485 3893 15519 3927
rect 15519 3893 15528 3927
rect 15476 3884 15528 3893
rect 16672 3927 16724 3936
rect 16672 3893 16681 3927
rect 16681 3893 16715 3927
rect 16715 3893 16724 3927
rect 16672 3884 16724 3893
rect 17224 3884 17276 3936
rect 17684 3884 17736 3936
rect 20352 4020 20404 4072
rect 21088 4097 21097 4131
rect 21097 4097 21131 4131
rect 21131 4097 21140 4131
rect 21088 4088 21140 4097
rect 24492 4088 24544 4140
rect 25964 4131 26016 4140
rect 25964 4097 25973 4131
rect 25973 4097 26007 4131
rect 26007 4097 26016 4131
rect 25964 4088 26016 4097
rect 27160 4088 27212 4140
rect 27344 4088 27396 4140
rect 30380 4156 30432 4208
rect 31208 4224 31260 4276
rect 32036 4224 32088 4276
rect 34336 4224 34388 4276
rect 34612 4224 34664 4276
rect 35072 4224 35124 4276
rect 35440 4224 35492 4276
rect 36544 4267 36596 4276
rect 36544 4233 36553 4267
rect 36553 4233 36587 4267
rect 36587 4233 36596 4267
rect 36544 4224 36596 4233
rect 21456 4020 21508 4072
rect 19616 3952 19668 4004
rect 20076 3952 20128 4004
rect 19524 3884 19576 3936
rect 21732 3952 21784 4004
rect 20352 3927 20404 3936
rect 20352 3893 20361 3927
rect 20361 3893 20395 3927
rect 20395 3893 20404 3927
rect 20352 3884 20404 3893
rect 20904 3927 20956 3936
rect 20904 3893 20913 3927
rect 20913 3893 20947 3927
rect 20947 3893 20956 3927
rect 20904 3884 20956 3893
rect 25688 4020 25740 4072
rect 24860 3952 24912 4004
rect 24952 3952 25004 4004
rect 22100 3884 22152 3936
rect 22560 3884 22612 3936
rect 25412 3884 25464 3936
rect 26424 3884 26476 3936
rect 27344 3952 27396 4004
rect 27528 3884 27580 3936
rect 27620 3884 27672 3936
rect 28356 3884 28408 3936
rect 31116 4156 31168 4208
rect 31668 4156 31720 4208
rect 36176 4156 36228 4208
rect 29460 4063 29512 4072
rect 29460 4029 29469 4063
rect 29469 4029 29503 4063
rect 29503 4029 29512 4063
rect 29460 4020 29512 4029
rect 29552 4020 29604 4072
rect 30748 4063 30800 4072
rect 30380 3952 30432 4004
rect 30748 4029 30757 4063
rect 30757 4029 30791 4063
rect 30791 4029 30800 4063
rect 30748 4020 30800 4029
rect 31208 4020 31260 4072
rect 31392 4088 31444 4140
rect 32312 4131 32364 4140
rect 32312 4097 32321 4131
rect 32321 4097 32355 4131
rect 32355 4097 32364 4131
rect 32312 4088 32364 4097
rect 34520 4131 34572 4140
rect 31668 4020 31720 4072
rect 29828 3927 29880 3936
rect 29828 3893 29837 3927
rect 29837 3893 29871 3927
rect 29871 3893 29880 3927
rect 29828 3884 29880 3893
rect 30472 3884 30524 3936
rect 34520 4097 34529 4131
rect 34529 4097 34563 4131
rect 34563 4097 34572 4131
rect 34520 4088 34572 4097
rect 34612 4088 34664 4140
rect 35808 4088 35860 4140
rect 36820 4088 36872 4140
rect 37648 4131 37700 4140
rect 37648 4097 37657 4131
rect 37657 4097 37691 4131
rect 37691 4097 37700 4131
rect 37648 4088 37700 4097
rect 33784 4020 33836 4072
rect 31484 3884 31536 3936
rect 32404 3884 32456 3936
rect 33876 3952 33928 4004
rect 35256 3952 35308 4004
rect 35624 3952 35676 4004
rect 32956 3884 33008 3936
rect 34796 3884 34848 3936
rect 37556 3884 37608 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 4620 3680 4672 3732
rect 8116 3680 8168 3732
rect 7564 3655 7616 3664
rect 7564 3621 7573 3655
rect 7573 3621 7607 3655
rect 7607 3621 7616 3655
rect 7564 3612 7616 3621
rect 1308 3476 1360 3528
rect 2412 3476 2464 3528
rect 3516 3476 3568 3528
rect 6460 3476 6512 3528
rect 7932 3476 7984 3528
rect 9588 3680 9640 3732
rect 11152 3723 11204 3732
rect 11152 3689 11161 3723
rect 11161 3689 11195 3723
rect 11195 3689 11204 3723
rect 11152 3680 11204 3689
rect 12532 3680 12584 3732
rect 14188 3680 14240 3732
rect 15660 3680 15712 3732
rect 16764 3680 16816 3732
rect 16948 3680 17000 3732
rect 19248 3680 19300 3732
rect 20720 3680 20772 3732
rect 21456 3680 21508 3732
rect 24584 3723 24636 3732
rect 8484 3612 8536 3664
rect 8944 3587 8996 3596
rect 8944 3553 8953 3587
rect 8953 3553 8987 3587
rect 8987 3553 8996 3587
rect 8944 3544 8996 3553
rect 9128 3587 9180 3596
rect 9128 3553 9137 3587
rect 9137 3553 9171 3587
rect 9171 3553 9180 3587
rect 9128 3544 9180 3553
rect 9634 3544 9686 3596
rect 17132 3612 17184 3664
rect 19892 3612 19944 3664
rect 24584 3689 24593 3723
rect 24593 3689 24627 3723
rect 24627 3689 24636 3723
rect 24584 3680 24636 3689
rect 26240 3680 26292 3732
rect 27160 3723 27212 3732
rect 27160 3689 27169 3723
rect 27169 3689 27203 3723
rect 27203 3689 27212 3723
rect 27160 3680 27212 3689
rect 27252 3680 27304 3732
rect 29920 3680 29972 3732
rect 30288 3680 30340 3732
rect 32312 3680 32364 3732
rect 32772 3680 32824 3732
rect 34060 3680 34112 3732
rect 12992 3544 13044 3596
rect 16948 3544 17000 3596
rect 17776 3544 17828 3596
rect 19064 3544 19116 3596
rect 19616 3544 19668 3596
rect 9036 3476 9088 3528
rect 9864 3476 9916 3528
rect 4620 3408 4672 3460
rect 9772 3408 9824 3460
rect 13544 3476 13596 3528
rect 14832 3476 14884 3528
rect 16856 3476 16908 3528
rect 2228 3340 2280 3392
rect 2872 3340 2924 3392
rect 8300 3383 8352 3392
rect 8300 3349 8309 3383
rect 8309 3349 8343 3383
rect 8343 3349 8352 3383
rect 8300 3340 8352 3349
rect 9680 3340 9732 3392
rect 12072 3408 12124 3460
rect 16672 3408 16724 3460
rect 9956 3340 10008 3392
rect 11060 3340 11112 3392
rect 13820 3340 13872 3392
rect 14648 3340 14700 3392
rect 15844 3340 15896 3392
rect 19432 3476 19484 3528
rect 22100 3544 22152 3596
rect 23572 3544 23624 3596
rect 29828 3612 29880 3664
rect 30564 3612 30616 3664
rect 30932 3612 30984 3664
rect 24952 3544 25004 3596
rect 23296 3476 23348 3528
rect 24400 3476 24452 3528
rect 25228 3476 25280 3528
rect 26700 3476 26752 3528
rect 27988 3519 28040 3528
rect 27988 3485 27997 3519
rect 27997 3485 28031 3519
rect 28031 3485 28040 3519
rect 27988 3476 28040 3485
rect 30012 3519 30064 3528
rect 30012 3485 30021 3519
rect 30021 3485 30055 3519
rect 30055 3485 30064 3519
rect 30012 3476 30064 3485
rect 30196 3476 30248 3528
rect 31024 3476 31076 3528
rect 31852 3519 31904 3528
rect 31852 3485 31861 3519
rect 31861 3485 31895 3519
rect 31895 3485 31904 3519
rect 31852 3476 31904 3485
rect 32036 3519 32088 3528
rect 32036 3485 32045 3519
rect 32045 3485 32079 3519
rect 32079 3485 32088 3519
rect 32036 3476 32088 3485
rect 32680 3544 32732 3596
rect 32220 3519 32272 3528
rect 32220 3485 32229 3519
rect 32229 3485 32263 3519
rect 32263 3485 32272 3519
rect 32220 3476 32272 3485
rect 32864 3476 32916 3528
rect 33048 3519 33100 3528
rect 33048 3485 33057 3519
rect 33057 3485 33091 3519
rect 33091 3485 33100 3519
rect 33048 3476 33100 3485
rect 33784 3519 33836 3528
rect 33784 3485 33793 3519
rect 33793 3485 33827 3519
rect 33827 3485 33836 3519
rect 33784 3476 33836 3485
rect 34428 3476 34480 3528
rect 34704 3519 34756 3528
rect 34704 3485 34713 3519
rect 34713 3485 34747 3519
rect 34747 3485 34756 3519
rect 34704 3476 34756 3485
rect 34796 3476 34848 3528
rect 35440 3476 35492 3528
rect 35716 3519 35768 3528
rect 35716 3485 35725 3519
rect 35725 3485 35759 3519
rect 35759 3485 35768 3519
rect 35716 3476 35768 3485
rect 36544 3519 36596 3528
rect 36544 3485 36553 3519
rect 36553 3485 36587 3519
rect 36587 3485 36596 3519
rect 36544 3476 36596 3485
rect 19524 3408 19576 3460
rect 20904 3408 20956 3460
rect 18328 3383 18380 3392
rect 18328 3349 18337 3383
rect 18337 3349 18371 3383
rect 18371 3349 18380 3383
rect 18328 3340 18380 3349
rect 19248 3340 19300 3392
rect 29828 3408 29880 3460
rect 28632 3383 28684 3392
rect 28632 3349 28641 3383
rect 28641 3349 28675 3383
rect 28675 3349 28684 3383
rect 28632 3340 28684 3349
rect 30840 3340 30892 3392
rect 32956 3408 33008 3460
rect 34336 3408 34388 3460
rect 35164 3408 35216 3460
rect 31116 3340 31168 3392
rect 32220 3340 32272 3392
rect 32312 3340 32364 3392
rect 35256 3340 35308 3392
rect 35440 3340 35492 3392
rect 36452 3340 36504 3392
rect 39396 3408 39448 3460
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 3056 3179 3108 3188
rect 3056 3145 3065 3179
rect 3065 3145 3099 3179
rect 3099 3145 3108 3179
rect 3056 3136 3108 3145
rect 4620 3179 4672 3188
rect 2872 3111 2924 3120
rect 2872 3077 2881 3111
rect 2881 3077 2915 3111
rect 2915 3077 2924 3111
rect 2872 3068 2924 3077
rect 4620 3145 4629 3179
rect 4629 3145 4663 3179
rect 4663 3145 4672 3179
rect 4620 3136 4672 3145
rect 5356 3136 5408 3188
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 3148 3000 3200 3052
rect 4620 3000 4672 3052
rect 6092 3000 6144 3052
rect 8760 3068 8812 3120
rect 8300 3000 8352 3052
rect 9128 3136 9180 3188
rect 9680 3136 9732 3188
rect 12348 3136 12400 3188
rect 12440 3136 12492 3188
rect 14280 3136 14332 3188
rect 9956 3000 10008 3052
rect 5540 2932 5592 2984
rect 11704 3111 11756 3120
rect 11704 3077 11713 3111
rect 11713 3077 11747 3111
rect 11747 3077 11756 3111
rect 11704 3068 11756 3077
rect 11796 3111 11848 3120
rect 11796 3077 11805 3111
rect 11805 3077 11839 3111
rect 11839 3077 11848 3111
rect 11796 3068 11848 3077
rect 2228 2864 2280 2916
rect 940 2796 992 2848
rect 2044 2796 2096 2848
rect 5356 2796 5408 2848
rect 11152 3000 11204 3052
rect 11888 3043 11940 3052
rect 11888 3009 11897 3043
rect 11897 3009 11931 3043
rect 11931 3009 11940 3043
rect 11888 3000 11940 3009
rect 12992 3068 13044 3120
rect 13360 3068 13412 3120
rect 14464 3068 14516 3120
rect 9680 2864 9732 2916
rect 10232 2864 10284 2916
rect 9864 2796 9916 2848
rect 10600 2796 10652 2848
rect 12716 3043 12768 3052
rect 12716 3009 12725 3043
rect 12725 3009 12759 3043
rect 12759 3009 12768 3043
rect 12716 3000 12768 3009
rect 13544 3000 13596 3052
rect 15200 3000 15252 3052
rect 16764 3000 16816 3052
rect 17684 3068 17736 3120
rect 18328 3068 18380 3120
rect 17868 3043 17920 3052
rect 12348 2932 12400 2984
rect 13268 2932 13320 2984
rect 14924 2864 14976 2916
rect 17868 3009 17877 3043
rect 17877 3009 17911 3043
rect 17911 3009 17920 3043
rect 17868 3000 17920 3009
rect 19156 3136 19208 3188
rect 22468 3136 22520 3188
rect 19984 3111 20036 3120
rect 19984 3077 19993 3111
rect 19993 3077 20027 3111
rect 20027 3077 20036 3111
rect 19984 3068 20036 3077
rect 20720 3043 20772 3052
rect 19248 2932 19300 2984
rect 20720 3009 20729 3043
rect 20729 3009 20763 3043
rect 20763 3009 20772 3043
rect 20720 3000 20772 3009
rect 20996 3043 21048 3052
rect 20996 3009 21005 3043
rect 21005 3009 21039 3043
rect 21039 3009 21048 3043
rect 20996 3000 21048 3009
rect 20352 2932 20404 2984
rect 12348 2796 12400 2848
rect 12624 2796 12676 2848
rect 14648 2796 14700 2848
rect 16856 2796 16908 2848
rect 21824 2864 21876 2916
rect 22376 3000 22428 3052
rect 23572 3043 23624 3052
rect 23572 3009 23581 3043
rect 23581 3009 23615 3043
rect 23615 3009 23624 3043
rect 23572 3000 23624 3009
rect 24952 3136 25004 3188
rect 25228 3136 25280 3188
rect 27896 3136 27948 3188
rect 28724 3179 28776 3188
rect 28724 3145 28733 3179
rect 28733 3145 28767 3179
rect 28767 3145 28776 3179
rect 28724 3136 28776 3145
rect 28816 3136 28868 3188
rect 35164 3136 35216 3188
rect 23848 3111 23900 3120
rect 23848 3077 23857 3111
rect 23857 3077 23891 3111
rect 23891 3077 23900 3111
rect 23848 3068 23900 3077
rect 19432 2796 19484 2848
rect 20812 2796 20864 2848
rect 23480 2796 23532 2848
rect 24860 3000 24912 3052
rect 25044 3043 25096 3052
rect 25044 3009 25053 3043
rect 25053 3009 25087 3043
rect 25087 3009 25096 3043
rect 25044 3000 25096 3009
rect 25320 3043 25372 3052
rect 25320 3009 25354 3043
rect 25354 3009 25372 3043
rect 25320 3000 25372 3009
rect 28632 3068 28684 3120
rect 30012 3068 30064 3120
rect 32036 3068 32088 3120
rect 29644 3043 29696 3052
rect 29644 3009 29653 3043
rect 29653 3009 29687 3043
rect 29687 3009 29696 3043
rect 29644 3000 29696 3009
rect 30932 3000 30984 3052
rect 31576 3000 31628 3052
rect 32864 3000 32916 3052
rect 35532 3000 35584 3052
rect 35256 2932 35308 2984
rect 38292 3000 38344 3052
rect 36912 2932 36964 2984
rect 25780 2796 25832 2848
rect 28080 2796 28132 2848
rect 31392 2864 31444 2916
rect 31024 2839 31076 2848
rect 31024 2805 31033 2839
rect 31033 2805 31067 2839
rect 31067 2805 31076 2839
rect 31024 2796 31076 2805
rect 31852 2796 31904 2848
rect 34704 2796 34756 2848
rect 35992 2839 36044 2848
rect 35992 2805 36001 2839
rect 36001 2805 36035 2839
rect 36035 2805 36044 2839
rect 35992 2796 36044 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 14832 2635 14884 2644
rect 1952 2499 2004 2508
rect 1952 2465 1961 2499
rect 1961 2465 1995 2499
rect 1995 2465 2004 2499
rect 1952 2456 2004 2465
rect 2780 2456 2832 2508
rect 12164 2524 12216 2576
rect 5264 2499 5316 2508
rect 5264 2465 5273 2499
rect 5273 2465 5307 2499
rect 5307 2465 5316 2499
rect 5264 2456 5316 2465
rect 4988 2431 5040 2440
rect 4988 2397 4997 2431
rect 4997 2397 5031 2431
rect 5031 2397 5040 2431
rect 4988 2388 5040 2397
rect 6920 2431 6972 2440
rect 6920 2397 6929 2431
rect 6929 2397 6963 2431
rect 6963 2397 6972 2431
rect 6920 2388 6972 2397
rect 7564 2388 7616 2440
rect 572 2320 624 2372
rect 11428 2456 11480 2508
rect 8944 2431 8996 2440
rect 8944 2397 8953 2431
rect 8953 2397 8987 2431
rect 8987 2397 8996 2431
rect 8944 2388 8996 2397
rect 10324 2388 10376 2440
rect 11520 2431 11572 2440
rect 3884 2252 3936 2304
rect 6828 2252 6880 2304
rect 9036 2320 9088 2372
rect 11520 2397 11529 2431
rect 11529 2397 11563 2431
rect 11563 2397 11572 2431
rect 11520 2388 11572 2397
rect 12992 2388 13044 2440
rect 14832 2601 14841 2635
rect 14841 2601 14875 2635
rect 14875 2601 14884 2635
rect 14832 2592 14884 2601
rect 17040 2635 17092 2644
rect 17040 2601 17049 2635
rect 17049 2601 17083 2635
rect 17083 2601 17092 2635
rect 17040 2592 17092 2601
rect 19524 2592 19576 2644
rect 21088 2592 21140 2644
rect 23296 2592 23348 2644
rect 25596 2592 25648 2644
rect 14188 2388 14240 2440
rect 14924 2456 14976 2508
rect 14464 2431 14516 2440
rect 14464 2397 14473 2431
rect 14473 2397 14507 2431
rect 14507 2397 14516 2431
rect 14464 2388 14516 2397
rect 14648 2431 14700 2440
rect 14648 2397 14657 2431
rect 14657 2397 14691 2431
rect 14691 2397 14700 2431
rect 14648 2388 14700 2397
rect 18880 2524 18932 2576
rect 20904 2524 20956 2576
rect 24308 2524 24360 2576
rect 24492 2499 24544 2508
rect 24492 2465 24501 2499
rect 24501 2465 24535 2499
rect 24535 2465 24544 2499
rect 24492 2456 24544 2465
rect 16856 2431 16908 2440
rect 16856 2397 16865 2431
rect 16865 2397 16899 2431
rect 16899 2397 16908 2431
rect 16856 2388 16908 2397
rect 18236 2388 18288 2440
rect 19432 2431 19484 2440
rect 8300 2252 8352 2304
rect 9772 2252 9824 2304
rect 10600 2295 10652 2304
rect 10600 2261 10609 2295
rect 10609 2261 10643 2295
rect 10643 2261 10652 2295
rect 10600 2252 10652 2261
rect 10876 2252 10928 2304
rect 11980 2252 12032 2304
rect 13084 2252 13136 2304
rect 15752 2320 15804 2372
rect 18144 2320 18196 2372
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 20812 2431 20864 2440
rect 20812 2397 20821 2431
rect 20821 2397 20855 2431
rect 20855 2397 20864 2431
rect 20812 2388 20864 2397
rect 20260 2320 20312 2372
rect 20444 2320 20496 2372
rect 21180 2320 21232 2372
rect 23480 2431 23532 2440
rect 23480 2397 23489 2431
rect 23489 2397 23523 2431
rect 23523 2397 23532 2431
rect 23480 2388 23532 2397
rect 25228 2388 25280 2440
rect 25780 2388 25832 2440
rect 27988 2592 28040 2644
rect 30196 2635 30248 2644
rect 30196 2601 30205 2635
rect 30205 2601 30239 2635
rect 30239 2601 30248 2635
rect 30196 2592 30248 2601
rect 30932 2592 30984 2644
rect 33048 2592 33100 2644
rect 27896 2431 27948 2440
rect 27896 2397 27905 2431
rect 27905 2397 27939 2431
rect 27939 2397 27948 2431
rect 27896 2388 27948 2397
rect 27988 2388 28040 2440
rect 28264 2431 28316 2440
rect 28264 2397 28273 2431
rect 28273 2397 28307 2431
rect 28307 2397 28316 2431
rect 28264 2388 28316 2397
rect 24860 2320 24912 2372
rect 25504 2363 25556 2372
rect 25504 2329 25513 2363
rect 25513 2329 25547 2363
rect 25547 2329 25556 2363
rect 25504 2320 25556 2329
rect 27344 2320 27396 2372
rect 29460 2320 29512 2372
rect 30380 2524 30432 2576
rect 31024 2524 31076 2576
rect 31116 2456 31168 2508
rect 32036 2456 32088 2508
rect 32956 2524 33008 2576
rect 33140 2524 33192 2576
rect 32220 2456 32272 2508
rect 30012 2431 30064 2440
rect 30012 2397 30021 2431
rect 30021 2397 30055 2431
rect 30055 2397 30064 2431
rect 30012 2388 30064 2397
rect 30656 2431 30708 2440
rect 30656 2397 30665 2431
rect 30665 2397 30699 2431
rect 30699 2397 30708 2431
rect 30656 2388 30708 2397
rect 30840 2388 30892 2440
rect 32312 2431 32364 2440
rect 32312 2397 32321 2431
rect 32321 2397 32355 2431
rect 32355 2397 32364 2431
rect 32312 2388 32364 2397
rect 33048 2456 33100 2508
rect 33692 2431 33744 2440
rect 33692 2397 33701 2431
rect 33701 2397 33735 2431
rect 33735 2397 33744 2431
rect 33692 2388 33744 2397
rect 33784 2388 33836 2440
rect 36084 2388 36136 2440
rect 36176 2431 36228 2440
rect 36176 2397 36185 2431
rect 36185 2397 36219 2431
rect 36219 2397 36228 2431
rect 36176 2388 36228 2397
rect 37188 2388 37240 2440
rect 31484 2320 31536 2372
rect 32036 2320 32088 2372
rect 16488 2252 16540 2304
rect 17592 2252 17644 2304
rect 18696 2252 18748 2304
rect 20076 2252 20128 2304
rect 24216 2252 24268 2304
rect 28724 2252 28776 2304
rect 30932 2252 30984 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 6920 2048 6972 2100
rect 10968 2048 11020 2100
rect 11520 2048 11572 2100
rect 16580 2048 16632 2100
rect 25504 2048 25556 2100
rect 27988 2048 28040 2100
rect 28172 2048 28224 2100
rect 33692 2048 33744 2100
rect 8944 1980 8996 2032
rect 15936 1980 15988 2032
rect 26608 1980 26660 2032
rect 33048 1980 33100 2032
rect 25780 1912 25832 1964
rect 28264 1912 28316 1964
rect 30012 1912 30064 1964
rect 24584 1368 24636 1420
rect 27436 1368 27488 1420
rect 34244 1368 34296 1420
rect 35992 1368 36044 1420
<< metal2 >>
rect 386 49200 442 50000
rect 1214 49200 1270 50000
rect 2042 49314 2098 50000
rect 2042 49286 2360 49314
rect 2042 49200 2098 49286
rect 400 47258 428 49200
rect 388 47252 440 47258
rect 388 47194 440 47200
rect 1228 46986 1256 49200
rect 2136 48204 2188 48210
rect 2136 48146 2188 48152
rect 1400 47660 1452 47666
rect 1400 47602 1452 47608
rect 1412 47054 1440 47602
rect 2148 47054 2176 48146
rect 2332 47258 2360 49286
rect 2870 49200 2926 50000
rect 3698 49314 3754 50000
rect 3698 49286 4016 49314
rect 3698 49200 3754 49286
rect 2320 47252 2372 47258
rect 2320 47194 2372 47200
rect 1400 47048 1452 47054
rect 1400 46990 1452 46996
rect 2136 47048 2188 47054
rect 2136 46990 2188 46996
rect 2884 47002 2912 49200
rect 3608 48136 3660 48142
rect 3608 48078 3660 48084
rect 3620 47054 3648 48078
rect 3792 48068 3844 48074
rect 3792 48010 3844 48016
rect 3804 47054 3832 48010
rect 3988 47190 4016 49286
rect 4526 49200 4582 50000
rect 5354 49200 5410 50000
rect 6182 49314 6238 50000
rect 7010 49314 7066 50000
rect 7838 49314 7894 50000
rect 6182 49286 6592 49314
rect 6182 49200 6238 49286
rect 4540 47546 4568 49200
rect 5080 47728 5132 47734
rect 5080 47670 5132 47676
rect 4540 47518 4660 47546
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4632 47258 4660 47518
rect 4620 47252 4672 47258
rect 4620 47194 4672 47200
rect 3976 47184 4028 47190
rect 3976 47126 4028 47132
rect 5092 47054 5120 47670
rect 5264 47524 5316 47530
rect 5264 47466 5316 47472
rect 5276 47054 5304 47466
rect 3608 47048 3660 47054
rect 2884 46986 3004 47002
rect 3608 46990 3660 46996
rect 3792 47048 3844 47054
rect 3792 46990 3844 46996
rect 5080 47048 5132 47054
rect 5080 46990 5132 46996
rect 5264 47048 5316 47054
rect 5264 46990 5316 46996
rect 1216 46980 1268 46986
rect 2884 46980 3016 46986
rect 2884 46974 2964 46980
rect 1216 46922 1268 46928
rect 2964 46922 3016 46928
rect 5368 46714 5396 49200
rect 6368 47796 6420 47802
rect 6368 47738 6420 47744
rect 6380 47054 6408 47738
rect 6564 47258 6592 49286
rect 7010 49286 7328 49314
rect 7010 49200 7066 49286
rect 7104 47456 7156 47462
rect 7104 47398 7156 47404
rect 6552 47252 6604 47258
rect 6552 47194 6604 47200
rect 7116 47054 7144 47398
rect 7300 47258 7328 49286
rect 7838 49286 8156 49314
rect 7838 49200 7894 49286
rect 8128 47258 8156 49286
rect 8666 49200 8722 50000
rect 9494 49314 9550 50000
rect 10322 49314 10378 50000
rect 9494 49286 9628 49314
rect 9494 49200 9550 49286
rect 8680 47258 8708 49200
rect 8944 47592 8996 47598
rect 8944 47534 8996 47540
rect 7288 47252 7340 47258
rect 7288 47194 7340 47200
rect 8116 47252 8168 47258
rect 8116 47194 8168 47200
rect 8668 47252 8720 47258
rect 8668 47194 8720 47200
rect 8956 47054 8984 47534
rect 9600 47240 9628 49286
rect 10322 49286 10640 49314
rect 10322 49200 10378 49286
rect 10416 47932 10468 47938
rect 10416 47874 10468 47880
rect 9680 47252 9732 47258
rect 9600 47212 9680 47240
rect 9680 47194 9732 47200
rect 10428 47054 10456 47874
rect 10612 47258 10640 49286
rect 11150 49200 11206 50000
rect 11978 49314 12034 50000
rect 11978 49286 12388 49314
rect 11978 49200 12034 49286
rect 11164 47258 11192 49200
rect 12072 47660 12124 47666
rect 12072 47602 12124 47608
rect 10600 47252 10652 47258
rect 10600 47194 10652 47200
rect 11152 47252 11204 47258
rect 11152 47194 11204 47200
rect 6368 47048 6420 47054
rect 6368 46990 6420 46996
rect 7104 47048 7156 47054
rect 7104 46990 7156 46996
rect 8944 47048 8996 47054
rect 8944 46990 8996 46996
rect 10416 47048 10468 47054
rect 10416 46990 10468 46996
rect 11520 47048 11572 47054
rect 11520 46990 11572 46996
rect 5356 46708 5408 46714
rect 5356 46650 5408 46656
rect 5448 46572 5500 46578
rect 5448 46514 5500 46520
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 5460 46170 5488 46514
rect 5448 46164 5500 46170
rect 5448 46106 5500 46112
rect 10692 46028 10744 46034
rect 10692 45970 10744 45976
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 10704 38010 10732 45970
rect 11532 41818 11560 46990
rect 11704 46504 11756 46510
rect 11704 46446 11756 46452
rect 11520 41812 11572 41818
rect 11520 41754 11572 41760
rect 11520 39976 11572 39982
rect 11520 39918 11572 39924
rect 11532 39098 11560 39918
rect 11612 39296 11664 39302
rect 11612 39238 11664 39244
rect 11520 39092 11572 39098
rect 11520 39034 11572 39040
rect 10692 38004 10744 38010
rect 10692 37946 10744 37952
rect 8944 37868 8996 37874
rect 8944 37810 8996 37816
rect 9588 37868 9640 37874
rect 9588 37810 9640 37816
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 8956 37330 8984 37810
rect 8944 37324 8996 37330
rect 8944 37266 8996 37272
rect 8956 36786 8984 37266
rect 9404 37188 9456 37194
rect 9404 37130 9456 37136
rect 8944 36780 8996 36786
rect 8944 36722 8996 36728
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 8944 34604 8996 34610
rect 8944 34546 8996 34552
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 5908 32428 5960 32434
rect 5908 32370 5960 32376
rect 8116 32428 8168 32434
rect 8116 32370 8168 32376
rect 5264 32224 5316 32230
rect 5264 32166 5316 32172
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4988 31816 5040 31822
rect 4988 31758 5040 31764
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 5000 30802 5028 31758
rect 5276 31754 5304 32166
rect 5264 31748 5316 31754
rect 5264 31690 5316 31696
rect 5920 31482 5948 32370
rect 6736 32360 6788 32366
rect 6736 32302 6788 32308
rect 6368 32224 6420 32230
rect 6368 32166 6420 32172
rect 6380 31754 6408 32166
rect 6288 31726 6408 31754
rect 5908 31476 5960 31482
rect 5908 31418 5960 31424
rect 5632 31136 5684 31142
rect 5632 31078 5684 31084
rect 5644 30938 5672 31078
rect 5632 30932 5684 30938
rect 5632 30874 5684 30880
rect 4988 30796 5040 30802
rect 4988 30738 5040 30744
rect 6288 30734 6316 31726
rect 6368 31680 6420 31686
rect 6368 31622 6420 31628
rect 6380 31142 6408 31622
rect 6748 31482 6776 32302
rect 7748 32224 7800 32230
rect 7748 32166 7800 32172
rect 7760 31822 7788 32166
rect 7012 31816 7064 31822
rect 7012 31758 7064 31764
rect 7748 31816 7800 31822
rect 7748 31758 7800 31764
rect 6828 31748 6880 31754
rect 6828 31690 6880 31696
rect 6552 31476 6604 31482
rect 6552 31418 6604 31424
rect 6736 31476 6788 31482
rect 6736 31418 6788 31424
rect 6368 31136 6420 31142
rect 6368 31078 6420 31084
rect 6276 30728 6328 30734
rect 6276 30670 6328 30676
rect 6368 30320 6420 30326
rect 6368 30262 6420 30268
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 5816 29844 5868 29850
rect 5816 29786 5868 29792
rect 5540 29572 5592 29578
rect 5540 29514 5592 29520
rect 4804 29504 4856 29510
rect 4804 29446 4856 29452
rect 5552 29458 5580 29514
rect 4816 29238 4844 29446
rect 5552 29430 5764 29458
rect 5540 29300 5592 29306
rect 5540 29242 5592 29248
rect 4804 29232 4856 29238
rect 4804 29174 4856 29180
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 5448 27464 5500 27470
rect 5552 27452 5580 29242
rect 5500 27424 5580 27452
rect 5448 27406 5500 27412
rect 5552 27062 5580 27424
rect 5540 27056 5592 27062
rect 5540 26998 5592 27004
rect 5448 26988 5500 26994
rect 5448 26930 5500 26936
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 5460 25498 5488 26930
rect 5552 26382 5580 26998
rect 5540 26376 5592 26382
rect 5540 26318 5592 26324
rect 5448 25492 5500 25498
rect 5448 25434 5500 25440
rect 4712 24812 4764 24818
rect 4712 24754 4764 24760
rect 4620 24608 4672 24614
rect 4620 24550 4672 24556
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4632 24138 4660 24550
rect 4620 24132 4672 24138
rect 4620 24074 4672 24080
rect 4724 23866 4752 24754
rect 5552 24274 5580 26318
rect 5632 26308 5684 26314
rect 5632 26250 5684 26256
rect 5644 26042 5672 26250
rect 5632 26036 5684 26042
rect 5632 25978 5684 25984
rect 5540 24268 5592 24274
rect 5540 24210 5592 24216
rect 5356 24064 5408 24070
rect 5356 24006 5408 24012
rect 4712 23860 4764 23866
rect 4712 23802 4764 23808
rect 4896 23724 4948 23730
rect 4896 23666 4948 23672
rect 4620 23520 4672 23526
rect 4620 23462 4672 23468
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4632 23118 4660 23462
rect 3792 23112 3844 23118
rect 3792 23054 3844 23060
rect 4620 23112 4672 23118
rect 4620 23054 4672 23060
rect 20 22568 72 22574
rect 20 22510 72 22516
rect 32 16574 60 22510
rect 3804 22030 3832 23054
rect 4712 22976 4764 22982
rect 4712 22918 4764 22924
rect 4724 22438 4752 22918
rect 4908 22506 4936 23666
rect 5368 23526 5396 24006
rect 5356 23520 5408 23526
rect 5356 23462 5408 23468
rect 5448 22704 5500 22710
rect 5448 22646 5500 22652
rect 4896 22500 4948 22506
rect 4896 22442 4948 22448
rect 4712 22432 4764 22438
rect 4712 22374 4764 22380
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 5460 22098 5488 22646
rect 5736 22642 5764 29430
rect 5828 29034 5856 29786
rect 5908 29504 5960 29510
rect 5908 29446 5960 29452
rect 5816 29028 5868 29034
rect 5816 28970 5868 28976
rect 5920 27470 5948 29446
rect 6380 29238 6408 30262
rect 6564 29238 6592 31418
rect 6736 31340 6788 31346
rect 6736 31282 6788 31288
rect 6748 30666 6776 31282
rect 6736 30660 6788 30666
rect 6736 30602 6788 30608
rect 6748 30326 6776 30602
rect 6736 30320 6788 30326
rect 6736 30262 6788 30268
rect 6736 29640 6788 29646
rect 6736 29582 6788 29588
rect 6368 29232 6420 29238
rect 6368 29174 6420 29180
rect 6552 29232 6604 29238
rect 6552 29174 6604 29180
rect 6380 28218 6408 29174
rect 6748 29034 6776 29582
rect 6840 29306 6868 31690
rect 7024 31346 7052 31758
rect 7012 31340 7064 31346
rect 7012 31282 7064 31288
rect 7288 31340 7340 31346
rect 7288 31282 7340 31288
rect 7300 30938 7328 31282
rect 8128 30938 8156 32370
rect 8956 31686 8984 34546
rect 9416 34202 9444 37130
rect 9600 34746 9628 37810
rect 10324 37120 10376 37126
rect 10322 37088 10324 37097
rect 10376 37088 10378 37097
rect 10322 37023 10378 37032
rect 9864 36780 9916 36786
rect 9864 36722 9916 36728
rect 9876 35290 9904 36722
rect 10336 35766 10364 37023
rect 10324 35760 10376 35766
rect 10324 35702 10376 35708
rect 9956 35488 10008 35494
rect 9956 35430 10008 35436
rect 9864 35284 9916 35290
rect 9864 35226 9916 35232
rect 9864 35148 9916 35154
rect 9864 35090 9916 35096
rect 9588 34740 9640 34746
rect 9588 34682 9640 34688
rect 9772 34536 9824 34542
rect 9772 34478 9824 34484
rect 9404 34196 9456 34202
rect 9404 34138 9456 34144
rect 9496 32836 9548 32842
rect 9496 32778 9548 32784
rect 9312 32360 9364 32366
rect 9312 32302 9364 32308
rect 9324 31822 9352 32302
rect 9508 32230 9536 32778
rect 9680 32768 9732 32774
rect 9680 32710 9732 32716
rect 9692 32502 9720 32710
rect 9680 32496 9732 32502
rect 9680 32438 9732 32444
rect 9496 32224 9548 32230
rect 9496 32166 9548 32172
rect 9036 31816 9088 31822
rect 9036 31758 9088 31764
rect 9312 31816 9364 31822
rect 9312 31758 9364 31764
rect 8392 31680 8444 31686
rect 8392 31622 8444 31628
rect 8944 31680 8996 31686
rect 8944 31622 8996 31628
rect 7288 30932 7340 30938
rect 7288 30874 7340 30880
rect 8116 30932 8168 30938
rect 8116 30874 8168 30880
rect 8404 30870 8432 31622
rect 8576 31136 8628 31142
rect 8576 31078 8628 31084
rect 8392 30864 8444 30870
rect 8392 30806 8444 30812
rect 7288 30728 7340 30734
rect 7288 30670 7340 30676
rect 7300 30394 7328 30670
rect 7932 30592 7984 30598
rect 7932 30534 7984 30540
rect 7288 30388 7340 30394
rect 7288 30330 7340 30336
rect 7944 30326 7972 30534
rect 7932 30320 7984 30326
rect 7932 30262 7984 30268
rect 8588 30122 8616 31078
rect 8576 30116 8628 30122
rect 8576 30058 8628 30064
rect 9048 29646 9076 31758
rect 9312 29708 9364 29714
rect 9312 29650 9364 29656
rect 8116 29640 8168 29646
rect 8116 29582 8168 29588
rect 9036 29640 9088 29646
rect 9036 29582 9088 29588
rect 7564 29504 7616 29510
rect 7564 29446 7616 29452
rect 6828 29300 6880 29306
rect 6828 29242 6880 29248
rect 6736 29028 6788 29034
rect 6736 28970 6788 28976
rect 6552 28960 6604 28966
rect 6552 28902 6604 28908
rect 6368 28212 6420 28218
rect 6368 28154 6420 28160
rect 6564 27674 6592 28902
rect 6840 28762 6868 29242
rect 6828 28756 6880 28762
rect 6828 28698 6880 28704
rect 7576 28082 7604 29446
rect 7932 29232 7984 29238
rect 7932 29174 7984 29180
rect 7944 28490 7972 29174
rect 8128 28694 8156 29582
rect 9048 29170 9076 29582
rect 9324 29578 9352 29650
rect 9312 29572 9364 29578
rect 9312 29514 9364 29520
rect 9036 29164 9088 29170
rect 9036 29106 9088 29112
rect 8668 28756 8720 28762
rect 8668 28698 8720 28704
rect 8116 28688 8168 28694
rect 8116 28630 8168 28636
rect 7748 28484 7800 28490
rect 7748 28426 7800 28432
rect 7932 28484 7984 28490
rect 7932 28426 7984 28432
rect 7196 28076 7248 28082
rect 7196 28018 7248 28024
rect 7564 28076 7616 28082
rect 7564 28018 7616 28024
rect 6552 27668 6604 27674
rect 6552 27610 6604 27616
rect 5908 27464 5960 27470
rect 5908 27406 5960 27412
rect 6920 27124 6972 27130
rect 6920 27066 6972 27072
rect 6460 27056 6512 27062
rect 6460 26998 6512 27004
rect 6472 25974 6500 26998
rect 6736 26784 6788 26790
rect 6736 26726 6788 26732
rect 6552 26240 6604 26246
rect 6552 26182 6604 26188
rect 6460 25968 6512 25974
rect 6460 25910 6512 25916
rect 6564 25702 6592 26182
rect 6552 25696 6604 25702
rect 6552 25638 6604 25644
rect 6748 25294 6776 26726
rect 6932 26042 6960 27066
rect 7208 26994 7236 28018
rect 7760 27402 7788 28426
rect 7944 27402 7972 28426
rect 8680 28218 8708 28698
rect 9048 28422 9076 29106
rect 9036 28416 9088 28422
rect 9036 28358 9088 28364
rect 8668 28212 8720 28218
rect 8668 28154 8720 28160
rect 9048 28082 9076 28358
rect 9036 28076 9088 28082
rect 9036 28018 9088 28024
rect 9220 28076 9272 28082
rect 9220 28018 9272 28024
rect 7748 27396 7800 27402
rect 7748 27338 7800 27344
rect 7932 27396 7984 27402
rect 7932 27338 7984 27344
rect 7760 27130 7788 27338
rect 8116 27328 8168 27334
rect 8116 27270 8168 27276
rect 7748 27124 7800 27130
rect 7748 27066 7800 27072
rect 8128 26994 8156 27270
rect 7196 26988 7248 26994
rect 7196 26930 7248 26936
rect 8116 26988 8168 26994
rect 8116 26930 8168 26936
rect 8668 26988 8720 26994
rect 8668 26930 8720 26936
rect 6920 26036 6972 26042
rect 6920 25978 6972 25984
rect 6736 25288 6788 25294
rect 6736 25230 6788 25236
rect 6644 25152 6696 25158
rect 6644 25094 6696 25100
rect 6184 24812 6236 24818
rect 6184 24754 6236 24760
rect 6196 24070 6224 24754
rect 6184 24064 6236 24070
rect 6184 24006 6236 24012
rect 6196 23798 6224 24006
rect 6184 23792 6236 23798
rect 6184 23734 6236 23740
rect 6656 23730 6684 25094
rect 6920 24880 6972 24886
rect 6920 24822 6972 24828
rect 6932 24138 6960 24822
rect 7104 24608 7156 24614
rect 7104 24550 7156 24556
rect 7116 24410 7144 24550
rect 7104 24404 7156 24410
rect 7104 24346 7156 24352
rect 6736 24132 6788 24138
rect 6736 24074 6788 24080
rect 6920 24132 6972 24138
rect 6920 24074 6972 24080
rect 6644 23724 6696 23730
rect 6644 23666 6696 23672
rect 6748 23322 6776 24074
rect 6932 23866 6960 24074
rect 6920 23860 6972 23866
rect 6920 23802 6972 23808
rect 6736 23316 6788 23322
rect 6736 23258 6788 23264
rect 7208 22642 7236 26930
rect 8484 26784 8536 26790
rect 8484 26726 8536 26732
rect 8496 26314 8524 26726
rect 8484 26308 8536 26314
rect 8484 26250 8536 26256
rect 8392 26240 8444 26246
rect 8392 26182 8444 26188
rect 8404 25770 8432 26182
rect 8680 26042 8708 26930
rect 9048 26382 9076 28018
rect 9232 27130 9260 28018
rect 9324 27334 9352 29514
rect 9508 28558 9536 32166
rect 9588 31748 9640 31754
rect 9588 31690 9640 31696
rect 9600 31482 9628 31690
rect 9588 31476 9640 31482
rect 9588 31418 9640 31424
rect 9680 31340 9732 31346
rect 9680 31282 9732 31288
rect 9692 30666 9720 31282
rect 9680 30660 9732 30666
rect 9680 30602 9732 30608
rect 9496 28552 9548 28558
rect 9496 28494 9548 28500
rect 9312 27328 9364 27334
rect 9312 27270 9364 27276
rect 9220 27124 9272 27130
rect 9220 27066 9272 27072
rect 9036 26376 9088 26382
rect 9036 26318 9088 26324
rect 8668 26036 8720 26042
rect 8668 25978 8720 25984
rect 9048 25906 9076 26318
rect 9036 25900 9088 25906
rect 9036 25842 9088 25848
rect 9588 25900 9640 25906
rect 9588 25842 9640 25848
rect 8392 25764 8444 25770
rect 8392 25706 8444 25712
rect 8392 25288 8444 25294
rect 8392 25230 8444 25236
rect 9036 25288 9088 25294
rect 9036 25230 9088 25236
rect 7288 24608 7340 24614
rect 7288 24550 7340 24556
rect 7300 23118 7328 24550
rect 8404 24410 8432 25230
rect 7748 24404 7800 24410
rect 7748 24346 7800 24352
rect 8392 24404 8444 24410
rect 8392 24346 8444 24352
rect 7380 24132 7432 24138
rect 7380 24074 7432 24080
rect 7288 23112 7340 23118
rect 7288 23054 7340 23060
rect 5724 22636 5776 22642
rect 5724 22578 5776 22584
rect 7196 22636 7248 22642
rect 7196 22578 7248 22584
rect 5448 22092 5500 22098
rect 5736 22094 5764 22578
rect 7012 22500 7064 22506
rect 7012 22442 7064 22448
rect 6920 22432 6972 22438
rect 6920 22374 6972 22380
rect 5736 22066 5856 22094
rect 5448 22034 5500 22040
rect 3792 22024 3844 22030
rect 3792 21966 3844 21972
rect 3804 20942 3832 21966
rect 5080 21548 5132 21554
rect 5080 21490 5132 21496
rect 4620 21344 4672 21350
rect 4620 21286 4672 21292
rect 4896 21344 4948 21350
rect 4896 21286 4948 21292
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 3792 20936 3844 20942
rect 3792 20878 3844 20884
rect 3804 20262 3832 20878
rect 4632 20534 4660 21286
rect 4908 20942 4936 21286
rect 4896 20936 4948 20942
rect 4896 20878 4948 20884
rect 4804 20800 4856 20806
rect 4804 20742 4856 20748
rect 4620 20528 4672 20534
rect 4620 20470 4672 20476
rect 2872 20256 2924 20262
rect 2872 20198 2924 20204
rect 3792 20256 3844 20262
rect 3792 20198 3844 20204
rect 2884 19922 2912 20198
rect 2872 19916 2924 19922
rect 2872 19858 2924 19864
rect 3804 19854 3832 20198
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 3792 19848 3844 19854
rect 3792 19790 3844 19796
rect 3804 18970 3832 19790
rect 4816 19174 4844 20742
rect 5092 19514 5120 21490
rect 5460 20618 5488 22034
rect 5724 21480 5776 21486
rect 5724 21422 5776 21428
rect 5368 20602 5580 20618
rect 5736 20602 5764 21422
rect 5368 20596 5592 20602
rect 5368 20590 5540 20596
rect 5080 19508 5132 19514
rect 5080 19450 5132 19456
rect 5368 19446 5396 20590
rect 5540 20538 5592 20544
rect 5724 20596 5776 20602
rect 5724 20538 5776 20544
rect 5448 20528 5500 20534
rect 5828 20482 5856 22066
rect 6276 21956 6328 21962
rect 6276 21898 6328 21904
rect 6288 21146 6316 21898
rect 6460 21480 6512 21486
rect 6460 21422 6512 21428
rect 6276 21140 6328 21146
rect 6276 21082 6328 21088
rect 6472 20534 6500 21422
rect 6932 20942 6960 22374
rect 7024 22234 7052 22442
rect 7012 22228 7064 22234
rect 7012 22170 7064 22176
rect 7208 22094 7236 22578
rect 7392 22506 7420 24074
rect 7760 23866 7788 24346
rect 9048 24070 9076 25230
rect 9600 24954 9628 25842
rect 9588 24948 9640 24954
rect 9588 24890 9640 24896
rect 9588 24404 9640 24410
rect 9588 24346 9640 24352
rect 8576 24064 8628 24070
rect 8576 24006 8628 24012
rect 9036 24064 9088 24070
rect 9036 24006 9088 24012
rect 9312 24064 9364 24070
rect 9312 24006 9364 24012
rect 7748 23860 7800 23866
rect 7748 23802 7800 23808
rect 8300 23724 8352 23730
rect 8300 23666 8352 23672
rect 8484 23724 8536 23730
rect 8484 23666 8536 23672
rect 8312 23186 8340 23666
rect 8496 23322 8524 23666
rect 8484 23316 8536 23322
rect 8484 23258 8536 23264
rect 8300 23180 8352 23186
rect 8300 23122 8352 23128
rect 7840 22704 7892 22710
rect 7840 22646 7892 22652
rect 7380 22500 7432 22506
rect 7380 22442 7432 22448
rect 7024 22066 7236 22094
rect 7024 21554 7052 22066
rect 7852 21690 7880 22646
rect 8588 22574 8616 24006
rect 9324 23202 9352 24006
rect 9600 23866 9628 24346
rect 9588 23860 9640 23866
rect 9588 23802 9640 23808
rect 8944 23180 8996 23186
rect 8944 23122 8996 23128
rect 9232 23174 9352 23202
rect 8668 22636 8720 22642
rect 8668 22578 8720 22584
rect 8576 22568 8628 22574
rect 8576 22510 8628 22516
rect 8680 22234 8708 22578
rect 8668 22228 8720 22234
rect 8668 22170 8720 22176
rect 8680 22098 8708 22170
rect 8668 22092 8720 22098
rect 8668 22034 8720 22040
rect 7564 21684 7616 21690
rect 7564 21626 7616 21632
rect 7840 21684 7892 21690
rect 7840 21626 7892 21632
rect 7380 21616 7432 21622
rect 7380 21558 7432 21564
rect 7012 21548 7064 21554
rect 7012 21490 7064 21496
rect 6920 20936 6972 20942
rect 6920 20878 6972 20884
rect 7024 20788 7052 21490
rect 7392 20874 7420 21558
rect 7380 20868 7432 20874
rect 7380 20810 7432 20816
rect 6932 20760 7052 20788
rect 5908 20528 5960 20534
rect 5500 20476 5908 20482
rect 5448 20470 5960 20476
rect 6460 20528 6512 20534
rect 6460 20470 6512 20476
rect 5460 20454 5948 20470
rect 5356 19440 5408 19446
rect 5356 19382 5408 19388
rect 5540 19440 5592 19446
rect 5540 19382 5592 19388
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 3792 18964 3844 18970
rect 3792 18906 3844 18912
rect 2688 17128 2740 17134
rect 2688 17070 2740 17076
rect 3700 17128 3752 17134
rect 3700 17070 3752 17076
rect 2700 16674 2728 17070
rect 2700 16658 2912 16674
rect 2700 16652 2924 16658
rect 2700 16646 2872 16652
rect 2700 16590 2728 16646
rect 2872 16594 2924 16600
rect 1860 16584 1912 16590
rect 32 16546 244 16574
rect 216 800 244 16546
rect 1860 16526 1912 16532
rect 2688 16584 2740 16590
rect 2688 16526 2740 16532
rect 1872 15570 1900 16526
rect 2700 16114 2728 16526
rect 2688 16108 2740 16114
rect 2688 16050 2740 16056
rect 1860 15564 1912 15570
rect 1860 15506 1912 15512
rect 2700 15026 2728 16050
rect 2688 15020 2740 15026
rect 2688 14962 2740 14968
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2700 13938 2728 14350
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2700 12850 2728 13874
rect 3712 12918 3740 17070
rect 3804 16658 3832 18906
rect 5368 18630 5396 19382
rect 5552 18970 5580 19382
rect 5644 19378 5672 20454
rect 6552 20256 6604 20262
rect 6552 20198 6604 20204
rect 6564 20058 6592 20198
rect 6552 20052 6604 20058
rect 6552 19994 6604 20000
rect 6932 19854 6960 20760
rect 7392 20534 7420 20810
rect 7576 20806 7604 21626
rect 8680 21554 8708 22034
rect 8668 21548 8720 21554
rect 8668 21490 8720 21496
rect 8956 21350 8984 23122
rect 9232 23118 9260 23174
rect 9220 23112 9272 23118
rect 9220 23054 9272 23060
rect 9692 22094 9720 30602
rect 9784 29714 9812 34478
rect 9876 34474 9904 35090
rect 9864 34468 9916 34474
rect 9864 34410 9916 34416
rect 9876 34134 9904 34410
rect 9864 34128 9916 34134
rect 9864 34070 9916 34076
rect 9876 33844 9904 34070
rect 9968 33998 9996 35430
rect 10508 35080 10560 35086
rect 10508 35022 10560 35028
rect 10416 34672 10468 34678
rect 10416 34614 10468 34620
rect 10232 34536 10284 34542
rect 10232 34478 10284 34484
rect 10244 33998 10272 34478
rect 9956 33992 10008 33998
rect 9956 33934 10008 33940
rect 10232 33992 10284 33998
rect 10232 33934 10284 33940
rect 9876 33816 9996 33844
rect 9968 33046 9996 33816
rect 9956 33040 10008 33046
rect 9956 32982 10008 32988
rect 9968 31482 9996 32982
rect 10244 32910 10272 33934
rect 10428 33658 10456 34614
rect 10520 34542 10548 35022
rect 10508 34536 10560 34542
rect 10508 34478 10560 34484
rect 10704 34354 10732 37946
rect 11624 37874 11652 39238
rect 11612 37868 11664 37874
rect 11612 37810 11664 37816
rect 11716 36582 11744 46446
rect 12084 45966 12112 47602
rect 12360 47240 12388 49286
rect 12806 49200 12862 50000
rect 13726 49200 13782 50000
rect 14554 49200 14610 50000
rect 15382 49200 15438 50000
rect 16210 49200 16266 50000
rect 17038 49200 17094 50000
rect 17866 49200 17922 50000
rect 18694 49200 18750 50000
rect 19522 49200 19578 50000
rect 20350 49314 20406 50000
rect 20350 49286 20668 49314
rect 20350 49200 20406 49286
rect 12716 47660 12768 47666
rect 12716 47602 12768 47608
rect 12440 47252 12492 47258
rect 12360 47212 12440 47240
rect 12440 47194 12492 47200
rect 12256 46572 12308 46578
rect 12256 46514 12308 46520
rect 12268 46170 12296 46514
rect 12256 46164 12308 46170
rect 12256 46106 12308 46112
rect 11980 45960 12032 45966
rect 11980 45902 12032 45908
rect 12072 45960 12124 45966
rect 12072 45902 12124 45908
rect 11888 38820 11940 38826
rect 11888 38762 11940 38768
rect 11796 38208 11848 38214
rect 11796 38150 11848 38156
rect 11152 36576 11204 36582
rect 11152 36518 11204 36524
rect 11704 36576 11756 36582
rect 11704 36518 11756 36524
rect 10968 35692 11020 35698
rect 10968 35634 11020 35640
rect 10980 35086 11008 35634
rect 11164 35193 11192 36518
rect 11612 36032 11664 36038
rect 11612 35974 11664 35980
rect 11624 35698 11652 35974
rect 11612 35692 11664 35698
rect 11612 35634 11664 35640
rect 11808 35290 11836 38150
rect 11900 37398 11928 38762
rect 11888 37392 11940 37398
rect 11888 37334 11940 37340
rect 11992 37346 12020 45902
rect 12084 40050 12112 45902
rect 12256 45484 12308 45490
rect 12256 45426 12308 45432
rect 12268 40730 12296 45426
rect 12256 40724 12308 40730
rect 12256 40666 12308 40672
rect 12532 40520 12584 40526
rect 12532 40462 12584 40468
rect 12072 40044 12124 40050
rect 12072 39986 12124 39992
rect 12544 39642 12572 40462
rect 12532 39636 12584 39642
rect 12532 39578 12584 39584
rect 12256 39432 12308 39438
rect 12256 39374 12308 39380
rect 12624 39432 12676 39438
rect 12624 39374 12676 39380
rect 11900 37210 11928 37334
rect 11992 37318 12112 37346
rect 11900 37182 12020 37210
rect 11888 37120 11940 37126
rect 11888 37062 11940 37068
rect 11900 36922 11928 37062
rect 11888 36916 11940 36922
rect 11888 36858 11940 36864
rect 11992 36650 12020 37182
rect 11980 36644 12032 36650
rect 11980 36586 12032 36592
rect 11796 35284 11848 35290
rect 11796 35226 11848 35232
rect 11150 35184 11206 35193
rect 11150 35119 11206 35128
rect 11164 35086 11192 35119
rect 10968 35080 11020 35086
rect 10968 35022 11020 35028
rect 11152 35080 11204 35086
rect 11152 35022 11204 35028
rect 10612 34326 10732 34354
rect 10416 33652 10468 33658
rect 10416 33594 10468 33600
rect 10612 33522 10640 34326
rect 10692 34196 10744 34202
rect 10692 34138 10744 34144
rect 10704 33998 10732 34138
rect 10980 34134 11008 35022
rect 12084 34728 12112 37318
rect 12268 37126 12296 39374
rect 12532 38888 12584 38894
rect 12532 38830 12584 38836
rect 12440 38412 12492 38418
rect 12440 38354 12492 38360
rect 12348 38004 12400 38010
rect 12348 37946 12400 37952
rect 12256 37120 12308 37126
rect 12256 37062 12308 37068
rect 12256 35488 12308 35494
rect 12256 35430 12308 35436
rect 12084 34700 12204 34728
rect 12072 34604 12124 34610
rect 12072 34546 12124 34552
rect 10968 34128 11020 34134
rect 10968 34070 11020 34076
rect 10692 33992 10744 33998
rect 10692 33934 10744 33940
rect 10600 33516 10652 33522
rect 10600 33458 10652 33464
rect 10232 32904 10284 32910
rect 10232 32846 10284 32852
rect 9956 31476 10008 31482
rect 9956 31418 10008 31424
rect 10244 31346 10272 32846
rect 10612 32842 10640 33458
rect 10600 32836 10652 32842
rect 10600 32778 10652 32784
rect 10232 31340 10284 31346
rect 10232 31282 10284 31288
rect 10232 30592 10284 30598
rect 10232 30534 10284 30540
rect 9772 29708 9824 29714
rect 9772 29650 9824 29656
rect 10244 29578 10272 30534
rect 10508 30252 10560 30258
rect 10508 30194 10560 30200
rect 10416 29844 10468 29850
rect 10416 29786 10468 29792
rect 10232 29572 10284 29578
rect 10232 29514 10284 29520
rect 10428 29306 10456 29786
rect 10416 29300 10468 29306
rect 10416 29242 10468 29248
rect 10520 29238 10548 30194
rect 10600 29504 10652 29510
rect 10600 29446 10652 29452
rect 10140 29232 10192 29238
rect 10140 29174 10192 29180
rect 10508 29232 10560 29238
rect 10508 29174 10560 29180
rect 9956 27464 10008 27470
rect 9956 27406 10008 27412
rect 9864 27396 9916 27402
rect 9864 27338 9916 27344
rect 9772 26784 9824 26790
rect 9772 26726 9824 26732
rect 9784 25974 9812 26726
rect 9772 25968 9824 25974
rect 9772 25910 9824 25916
rect 9784 25158 9812 25910
rect 9876 25498 9904 27338
rect 9968 26994 9996 27406
rect 9956 26988 10008 26994
rect 9956 26930 10008 26936
rect 9864 25492 9916 25498
rect 9864 25434 9916 25440
rect 9772 25152 9824 25158
rect 9772 25094 9824 25100
rect 9968 24410 9996 26930
rect 10048 26240 10100 26246
rect 10048 26182 10100 26188
rect 10060 25498 10088 26182
rect 10048 25492 10100 25498
rect 10048 25434 10100 25440
rect 9956 24404 10008 24410
rect 9956 24346 10008 24352
rect 10152 24342 10180 29174
rect 10416 29164 10468 29170
rect 10416 29106 10468 29112
rect 10428 27130 10456 29106
rect 10508 27872 10560 27878
rect 10508 27814 10560 27820
rect 10520 27674 10548 27814
rect 10508 27668 10560 27674
rect 10508 27610 10560 27616
rect 10416 27124 10468 27130
rect 10416 27066 10468 27072
rect 10612 26994 10640 29446
rect 10600 26988 10652 26994
rect 10600 26930 10652 26936
rect 10232 25900 10284 25906
rect 10232 25842 10284 25848
rect 10244 25498 10272 25842
rect 10324 25696 10376 25702
rect 10324 25638 10376 25644
rect 10336 25498 10364 25638
rect 10232 25492 10284 25498
rect 10232 25434 10284 25440
rect 10324 25492 10376 25498
rect 10324 25434 10376 25440
rect 10140 24336 10192 24342
rect 10140 24278 10192 24284
rect 10152 24070 10180 24278
rect 10140 24064 10192 24070
rect 10140 24006 10192 24012
rect 10600 23520 10652 23526
rect 10600 23462 10652 23468
rect 10612 23322 10640 23462
rect 10600 23316 10652 23322
rect 10600 23258 10652 23264
rect 10048 23044 10100 23050
rect 10048 22986 10100 22992
rect 10060 22506 10088 22986
rect 10048 22500 10100 22506
rect 10048 22442 10100 22448
rect 10704 22094 10732 33934
rect 10980 33590 11008 34070
rect 11980 33992 12032 33998
rect 11980 33934 12032 33940
rect 11520 33924 11572 33930
rect 11520 33866 11572 33872
rect 10784 33584 10836 33590
rect 10784 33526 10836 33532
rect 10968 33584 11020 33590
rect 10968 33526 11020 33532
rect 11060 33584 11112 33590
rect 11060 33526 11112 33532
rect 10796 32910 10824 33526
rect 11072 32910 11100 33526
rect 10784 32904 10836 32910
rect 10784 32846 10836 32852
rect 11060 32904 11112 32910
rect 11060 32846 11112 32852
rect 10796 32502 10824 32846
rect 11072 32570 11100 32846
rect 11060 32564 11112 32570
rect 11060 32506 11112 32512
rect 10784 32496 10836 32502
rect 10784 32438 10836 32444
rect 11060 32224 11112 32230
rect 11060 32166 11112 32172
rect 11072 31278 11100 32166
rect 11532 31754 11560 33866
rect 11992 33658 12020 33934
rect 11980 33652 12032 33658
rect 11980 33594 12032 33600
rect 12084 33046 12112 34546
rect 12176 33658 12204 34700
rect 12268 34610 12296 35430
rect 12256 34604 12308 34610
rect 12256 34546 12308 34552
rect 12360 33998 12388 37946
rect 12452 37942 12480 38354
rect 12544 38214 12572 38830
rect 12532 38208 12584 38214
rect 12532 38150 12584 38156
rect 12440 37936 12492 37942
rect 12440 37878 12492 37884
rect 12452 35766 12480 37878
rect 12532 36780 12584 36786
rect 12532 36722 12584 36728
rect 12440 35760 12492 35766
rect 12544 35737 12572 36722
rect 12440 35702 12492 35708
rect 12530 35728 12586 35737
rect 12530 35663 12586 35672
rect 12440 35012 12492 35018
rect 12440 34954 12492 34960
rect 12348 33992 12400 33998
rect 12348 33934 12400 33940
rect 12164 33652 12216 33658
rect 12164 33594 12216 33600
rect 12452 33590 12480 34954
rect 12636 34746 12664 39374
rect 12728 38554 12756 47602
rect 12820 47258 12848 49200
rect 13176 48136 13228 48142
rect 13176 48078 13228 48084
rect 12992 48000 13044 48006
rect 12992 47942 13044 47948
rect 12808 47252 12860 47258
rect 12808 47194 12860 47200
rect 13004 47054 13032 47942
rect 12992 47048 13044 47054
rect 12992 46990 13044 46996
rect 13188 45948 13216 48078
rect 13740 47240 13768 49200
rect 14004 48204 14056 48210
rect 14004 48146 14056 48152
rect 13912 47456 13964 47462
rect 13912 47398 13964 47404
rect 13820 47252 13872 47258
rect 13740 47212 13820 47240
rect 13820 47194 13872 47200
rect 13268 47048 13320 47054
rect 13268 46990 13320 46996
rect 13280 46714 13308 46990
rect 13268 46708 13320 46714
rect 13268 46650 13320 46656
rect 13268 45960 13320 45966
rect 13188 45920 13268 45948
rect 13268 45902 13320 45908
rect 13280 45626 13308 45902
rect 13924 45898 13952 47398
rect 14016 46578 14044 48146
rect 14568 47258 14596 49200
rect 15108 48068 15160 48074
rect 15108 48010 15160 48016
rect 14556 47252 14608 47258
rect 14556 47194 14608 47200
rect 14832 47048 14884 47054
rect 14832 46990 14884 46996
rect 14004 46572 14056 46578
rect 14004 46514 14056 46520
rect 14464 46572 14516 46578
rect 14464 46514 14516 46520
rect 13912 45892 13964 45898
rect 13912 45834 13964 45840
rect 13268 45620 13320 45626
rect 13268 45562 13320 45568
rect 13544 45416 13596 45422
rect 13544 45358 13596 45364
rect 12900 44328 12952 44334
rect 12900 44270 12952 44276
rect 12912 40050 12940 44270
rect 13268 42628 13320 42634
rect 13268 42570 13320 42576
rect 13280 41478 13308 42570
rect 13268 41472 13320 41478
rect 13268 41414 13320 41420
rect 13452 41472 13504 41478
rect 13452 41414 13504 41420
rect 13280 41274 13308 41414
rect 13372 41386 13492 41414
rect 13268 41268 13320 41274
rect 13268 41210 13320 41216
rect 13176 41200 13228 41206
rect 13176 41142 13228 41148
rect 12992 41064 13044 41070
rect 12992 41006 13044 41012
rect 12900 40044 12952 40050
rect 12900 39986 12952 39992
rect 12716 38548 12768 38554
rect 12716 38490 12768 38496
rect 12912 38418 12940 39986
rect 12900 38412 12952 38418
rect 12900 38354 12952 38360
rect 12716 38276 12768 38282
rect 12716 38218 12768 38224
rect 12728 35222 12756 38218
rect 12808 36712 12860 36718
rect 12808 36654 12860 36660
rect 12716 35216 12768 35222
rect 12716 35158 12768 35164
rect 12624 34740 12676 34746
rect 12624 34682 12676 34688
rect 12624 34604 12676 34610
rect 12624 34546 12676 34552
rect 12636 33998 12664 34546
rect 12624 33992 12676 33998
rect 12624 33934 12676 33940
rect 12624 33856 12676 33862
rect 12624 33798 12676 33804
rect 12440 33584 12492 33590
rect 12440 33526 12492 33532
rect 12164 33516 12216 33522
rect 12164 33458 12216 33464
rect 12072 33040 12124 33046
rect 12072 32982 12124 32988
rect 12176 32978 12204 33458
rect 12348 33448 12400 33454
rect 12348 33390 12400 33396
rect 12360 33289 12388 33390
rect 12346 33280 12402 33289
rect 12346 33215 12402 33224
rect 12164 32972 12216 32978
rect 12164 32914 12216 32920
rect 12360 32910 12388 33215
rect 12348 32904 12400 32910
rect 12348 32846 12400 32852
rect 11888 32768 11940 32774
rect 11888 32710 11940 32716
rect 11704 32428 11756 32434
rect 11704 32370 11756 32376
rect 11716 32026 11744 32370
rect 11704 32020 11756 32026
rect 11704 31962 11756 31968
rect 11440 31726 11560 31754
rect 11060 31272 11112 31278
rect 11060 31214 11112 31220
rect 10876 30320 10928 30326
rect 10876 30262 10928 30268
rect 10888 29646 10916 30262
rect 10876 29640 10928 29646
rect 10876 29582 10928 29588
rect 10784 28212 10836 28218
rect 10784 28154 10836 28160
rect 10796 27470 10824 28154
rect 10888 27606 10916 29582
rect 10876 27600 10928 27606
rect 10876 27542 10928 27548
rect 11440 27470 11468 31726
rect 11796 29844 11848 29850
rect 11796 29786 11848 29792
rect 11612 29572 11664 29578
rect 11612 29514 11664 29520
rect 11624 29306 11652 29514
rect 11612 29300 11664 29306
rect 11612 29242 11664 29248
rect 11808 29170 11836 29786
rect 11900 29578 11928 32710
rect 11980 32360 12032 32366
rect 11980 32302 12032 32308
rect 11992 32026 12020 32302
rect 11980 32020 12032 32026
rect 11980 31962 12032 31968
rect 11992 30802 12020 31962
rect 11980 30796 12032 30802
rect 11980 30738 12032 30744
rect 11888 29572 11940 29578
rect 11888 29514 11940 29520
rect 11900 29306 11928 29514
rect 11888 29300 11940 29306
rect 11888 29242 11940 29248
rect 11796 29164 11848 29170
rect 11796 29106 11848 29112
rect 11888 28960 11940 28966
rect 11888 28902 11940 28908
rect 11520 28416 11572 28422
rect 11520 28358 11572 28364
rect 11532 28082 11560 28358
rect 11520 28076 11572 28082
rect 11520 28018 11572 28024
rect 11612 28076 11664 28082
rect 11612 28018 11664 28024
rect 10784 27464 10836 27470
rect 10784 27406 10836 27412
rect 11428 27464 11480 27470
rect 11428 27406 11480 27412
rect 10784 26308 10836 26314
rect 10784 26250 10836 26256
rect 10796 26042 10824 26250
rect 10784 26036 10836 26042
rect 10784 25978 10836 25984
rect 10784 25220 10836 25226
rect 10784 25162 10836 25168
rect 10796 23866 10824 25162
rect 11060 25152 11112 25158
rect 11060 25094 11112 25100
rect 11072 24886 11100 25094
rect 11060 24880 11112 24886
rect 11060 24822 11112 24828
rect 10784 23860 10836 23866
rect 10784 23802 10836 23808
rect 11440 23730 11468 27406
rect 11532 26586 11560 28018
rect 11624 27674 11652 28018
rect 11612 27668 11664 27674
rect 11612 27610 11664 27616
rect 11900 27470 11928 28902
rect 11888 27464 11940 27470
rect 11888 27406 11940 27412
rect 11520 26580 11572 26586
rect 11520 26522 11572 26528
rect 11992 25294 12020 30738
rect 12452 29850 12480 33526
rect 12532 30388 12584 30394
rect 12532 30330 12584 30336
rect 12440 29844 12492 29850
rect 12440 29786 12492 29792
rect 12072 29504 12124 29510
rect 12072 29446 12124 29452
rect 12084 29170 12112 29446
rect 12176 29294 12480 29322
rect 12072 29164 12124 29170
rect 12072 29106 12124 29112
rect 12176 28422 12204 29294
rect 12452 29238 12480 29294
rect 12348 29232 12400 29238
rect 12346 29200 12348 29209
rect 12440 29232 12492 29238
rect 12400 29200 12402 29209
rect 12440 29174 12492 29180
rect 12346 29135 12402 29144
rect 12544 29050 12572 30330
rect 12452 29022 12572 29050
rect 12452 28994 12480 29022
rect 12360 28966 12480 28994
rect 12164 28416 12216 28422
rect 12164 28358 12216 28364
rect 11980 25288 12032 25294
rect 11980 25230 12032 25236
rect 11704 25152 11756 25158
rect 11704 25094 11756 25100
rect 12164 25152 12216 25158
rect 12164 25094 12216 25100
rect 11520 24200 11572 24206
rect 11520 24142 11572 24148
rect 11532 23866 11560 24142
rect 11520 23860 11572 23866
rect 11520 23802 11572 23808
rect 11428 23724 11480 23730
rect 11428 23666 11480 23672
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 10796 22642 10824 23462
rect 10784 22636 10836 22642
rect 10784 22578 10836 22584
rect 11244 22636 11296 22642
rect 11244 22578 11296 22584
rect 9692 22066 9904 22094
rect 9220 21548 9272 21554
rect 9220 21490 9272 21496
rect 8300 21344 8352 21350
rect 8300 21286 8352 21292
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 7564 20800 7616 20806
rect 7564 20742 7616 20748
rect 7576 20534 7604 20742
rect 7380 20528 7432 20534
rect 7380 20470 7432 20476
rect 7564 20528 7616 20534
rect 7564 20470 7616 20476
rect 6920 19848 6972 19854
rect 6920 19790 6972 19796
rect 6460 19712 6512 19718
rect 6460 19654 6512 19660
rect 5632 19372 5684 19378
rect 5632 19314 5684 19320
rect 5816 19372 5868 19378
rect 5816 19314 5868 19320
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5828 18902 5856 19314
rect 5816 18896 5868 18902
rect 5816 18838 5868 18844
rect 6472 18698 6500 19654
rect 6460 18692 6512 18698
rect 6460 18634 6512 18640
rect 5356 18624 5408 18630
rect 5356 18566 5408 18572
rect 6932 18426 6960 19790
rect 7392 19786 7420 20470
rect 7576 19786 7604 20470
rect 7380 19780 7432 19786
rect 7380 19722 7432 19728
rect 7564 19780 7616 19786
rect 7564 19722 7616 19728
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7760 18970 7788 19110
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 8312 18766 8340 21286
rect 8956 21010 8984 21286
rect 8944 21004 8996 21010
rect 8944 20946 8996 20952
rect 8484 20936 8536 20942
rect 8484 20878 8536 20884
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 8404 19854 8432 20198
rect 8496 19990 8524 20878
rect 8956 20534 8984 20946
rect 9036 20800 9088 20806
rect 9036 20742 9088 20748
rect 8944 20528 8996 20534
rect 8944 20470 8996 20476
rect 8668 20460 8720 20466
rect 8668 20402 8720 20408
rect 8680 20058 8708 20402
rect 8668 20052 8720 20058
rect 8668 19994 8720 20000
rect 8484 19984 8536 19990
rect 8484 19926 8536 19932
rect 8956 19922 8984 20470
rect 8944 19916 8996 19922
rect 8944 19858 8996 19864
rect 8392 19848 8444 19854
rect 8392 19790 8444 19796
rect 8956 19446 8984 19858
rect 9048 19854 9076 20742
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 9232 19446 9260 21490
rect 9496 21412 9548 21418
rect 9496 21354 9548 21360
rect 9508 19514 9536 21354
rect 9588 21140 9640 21146
rect 9588 21082 9640 21088
rect 9600 20466 9628 21082
rect 9588 20460 9640 20466
rect 9588 20402 9640 20408
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 8944 19440 8996 19446
rect 8944 19382 8996 19388
rect 9220 19440 9272 19446
rect 9220 19382 9272 19388
rect 8668 19372 8720 19378
rect 8668 19314 8720 19320
rect 8680 18970 8708 19314
rect 8668 18964 8720 18970
rect 8668 18906 8720 18912
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 5908 17808 5960 17814
rect 5908 17750 5960 17756
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 3792 16652 3844 16658
rect 3792 16594 3844 16600
rect 4080 16590 4108 17274
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 4620 17060 4672 17066
rect 4620 17002 4672 17008
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3804 14482 3832 15438
rect 3884 15428 3936 15434
rect 3884 15370 3936 15376
rect 3896 15162 3924 15370
rect 3884 15156 3936 15162
rect 3884 15098 3936 15104
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 4632 14414 4660 17002
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 4724 14618 4752 16118
rect 5092 15978 5120 16390
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 5080 15972 5132 15978
rect 5080 15914 5132 15920
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 5262 15872 5318 15881
rect 4816 15434 4844 15846
rect 5262 15807 5318 15816
rect 4804 15428 4856 15434
rect 4804 15370 4856 15376
rect 4804 14884 4856 14890
rect 4804 14826 4856 14832
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4816 14006 4844 14826
rect 5276 14226 5304 15807
rect 5368 15026 5396 16050
rect 5356 15020 5408 15026
rect 5356 14962 5408 14968
rect 5368 14550 5396 14962
rect 5356 14544 5408 14550
rect 5356 14486 5408 14492
rect 5276 14198 5396 14226
rect 4804 14000 4856 14006
rect 4804 13942 4856 13948
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 3700 12912 3752 12918
rect 3700 12854 3752 12860
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 1400 9920 1452 9926
rect 1400 9862 1452 9868
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 940 2848 992 2854
rect 940 2790 992 2796
rect 572 2372 624 2378
rect 572 2314 624 2320
rect 584 800 612 2314
rect 952 800 980 2790
rect 1320 800 1348 3470
rect 1412 3058 1440 9862
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1688 800 1716 3878
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2240 2922 2268 3334
rect 2228 2916 2280 2922
rect 2228 2858 2280 2864
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 1950 2544 2006 2553
rect 1950 2479 1952 2488
rect 2004 2479 2006 2488
rect 1952 2450 2004 2456
rect 2056 800 2084 2790
rect 2424 800 2452 3470
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 2884 3126 2912 3334
rect 3068 3194 3096 3878
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4632 3738 4660 8502
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 2872 3120 2924 3126
rect 2872 3062 2924 3068
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2792 800 2820 2450
rect 3160 800 3188 2994
rect 3528 800 3556 3470
rect 4620 3460 4672 3466
rect 4620 3402 4672 3408
rect 4632 3194 4660 3402
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 3896 800 3924 2246
rect 4632 800 4660 2994
rect 5276 2514 5304 12718
rect 5368 3194 5396 14198
rect 5460 13530 5488 17138
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5552 15026 5580 16934
rect 5724 16516 5776 16522
rect 5724 16458 5776 16464
rect 5632 16448 5684 16454
rect 5632 16390 5684 16396
rect 5540 15020 5592 15026
rect 5540 14962 5592 14968
rect 5644 14074 5672 16390
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 5736 13870 5764 16458
rect 5828 16182 5856 17614
rect 5816 16176 5868 16182
rect 5816 16118 5868 16124
rect 5920 15434 5948 17750
rect 7104 17672 7156 17678
rect 7104 17614 7156 17620
rect 6184 17536 6236 17542
rect 6184 17478 6236 17484
rect 6092 17264 6144 17270
rect 6092 17206 6144 17212
rect 6000 16516 6052 16522
rect 6000 16458 6052 16464
rect 6012 16114 6040 16458
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 5908 15428 5960 15434
rect 5908 15370 5960 15376
rect 6000 15428 6052 15434
rect 6000 15370 6052 15376
rect 6012 15094 6040 15370
rect 6000 15088 6052 15094
rect 6000 15030 6052 15036
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 6104 12986 6132 17206
rect 6196 14482 6224 17478
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 7024 16522 7052 17138
rect 7012 16516 7064 16522
rect 7012 16458 7064 16464
rect 6368 16108 6420 16114
rect 6368 16050 6420 16056
rect 6276 16040 6328 16046
rect 6276 15982 6328 15988
rect 6184 14476 6236 14482
rect 6184 14418 6236 14424
rect 6288 14074 6316 15982
rect 6380 15026 6408 16050
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6644 15972 6696 15978
rect 6644 15914 6696 15920
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6368 15020 6420 15026
rect 6368 14962 6420 14968
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 6380 13938 6408 14962
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6472 13326 6500 14758
rect 6564 13938 6592 15302
rect 6656 14958 6684 15914
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 6644 14952 6696 14958
rect 6644 14894 6696 14900
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 6656 14006 6684 14758
rect 6644 14000 6696 14006
rect 6644 13942 6696 13948
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6748 13870 6776 15506
rect 6840 15502 6868 15982
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6828 15496 6880 15502
rect 6828 15438 6880 15444
rect 6840 14278 6868 15438
rect 6932 15094 6960 15846
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6840 13326 6868 14214
rect 7024 14006 7052 15302
rect 7116 14074 7144 17614
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7392 16794 7420 17138
rect 8116 17128 8168 17134
rect 8116 17070 8168 17076
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 7012 14000 7064 14006
rect 7012 13942 7064 13948
rect 7208 13938 7236 16390
rect 7840 16244 7892 16250
rect 7840 16186 7892 16192
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 7288 15904 7340 15910
rect 7286 15872 7288 15881
rect 7340 15872 7342 15881
rect 7286 15807 7342 15816
rect 7392 15162 7420 16050
rect 7380 15156 7432 15162
rect 7380 15098 7432 15104
rect 7852 15026 7880 16186
rect 8024 16176 8076 16182
rect 8024 16118 8076 16124
rect 8036 15162 8064 16118
rect 8024 15156 8076 15162
rect 8024 15098 8076 15104
rect 7840 15020 7892 15026
rect 7840 14962 7892 14968
rect 7932 14952 7984 14958
rect 7852 14900 7932 14906
rect 7852 14894 7984 14900
rect 7852 14878 7972 14894
rect 7852 14346 7880 14878
rect 8128 14618 8156 17070
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 8220 16182 8248 16934
rect 8208 16176 8260 16182
rect 8208 16118 8260 16124
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8220 14822 8248 15098
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8116 14612 8168 14618
rect 8116 14554 8168 14560
rect 8220 14482 8248 14758
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 7840 14340 7892 14346
rect 7840 14282 7892 14288
rect 7852 13938 7880 14282
rect 8116 14000 8168 14006
rect 8116 13942 8168 13948
rect 7196 13932 7248 13938
rect 7196 13874 7248 13880
rect 7840 13932 7892 13938
rect 7840 13874 7892 13880
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6840 12850 6868 13262
rect 7932 13252 7984 13258
rect 7932 13194 7984 13200
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6840 12306 6868 12786
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 7944 11898 7972 13194
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 8128 11762 8156 13942
rect 8220 13938 8248 14418
rect 8404 14414 8432 18770
rect 8956 18290 8984 19382
rect 9232 18834 9260 19382
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 8864 17882 8892 18226
rect 8852 17876 8904 17882
rect 8852 17818 8904 17824
rect 8864 17134 8892 17818
rect 9404 17808 9456 17814
rect 9404 17750 9456 17756
rect 9416 17610 9444 17750
rect 9404 17604 9456 17610
rect 9404 17546 9456 17552
rect 9416 17513 9444 17546
rect 9402 17504 9458 17513
rect 9402 17439 9458 17448
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8864 16726 8892 17070
rect 9324 16794 9352 17138
rect 9036 16788 9088 16794
rect 9036 16730 9088 16736
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 8852 16720 8904 16726
rect 8852 16662 8904 16668
rect 8944 16516 8996 16522
rect 8944 16458 8996 16464
rect 8956 15502 8984 16458
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 8852 15360 8904 15366
rect 8852 15302 8904 15308
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8312 12442 8340 13874
rect 8404 12986 8432 14350
rect 8864 13258 8892 15302
rect 8956 15026 8984 15438
rect 9048 15026 9076 16730
rect 9128 16516 9180 16522
rect 9128 16458 9180 16464
rect 9140 16250 9168 16458
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 9416 16250 9444 16390
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9784 15502 9812 15642
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 8944 15020 8996 15026
rect 8944 14962 8996 14968
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 9784 14482 9812 15438
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8852 13252 8904 13258
rect 8852 13194 8904 13200
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8956 12918 8984 14214
rect 9140 13530 9168 14350
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9232 13462 9260 13874
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9220 13456 9272 13462
rect 9220 13398 9272 13404
rect 9128 13252 9180 13258
rect 9128 13194 9180 13200
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 8944 12912 8996 12918
rect 8944 12854 8996 12860
rect 8300 12436 8352 12442
rect 9048 12434 9076 12922
rect 9140 12714 9168 13194
rect 9128 12708 9180 12714
rect 9128 12650 9180 12656
rect 9048 12406 9260 12434
rect 8300 12378 8352 12384
rect 9232 11830 9260 12406
rect 9784 12238 9812 13806
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9220 11824 9272 11830
rect 9220 11766 9272 11772
rect 8116 11756 8168 11762
rect 8116 11698 8168 11704
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7484 7818 7512 8230
rect 7472 7812 7524 7818
rect 7472 7754 7524 7760
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5552 2990 5580 5646
rect 7576 3670 7604 10746
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 8956 9654 8984 9862
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 7932 9512 7984 9518
rect 9048 9466 9076 9862
rect 7932 9454 7984 9460
rect 7944 9042 7972 9454
rect 8864 9438 9076 9466
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 7944 7886 7972 8978
rect 8220 8498 8248 9318
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8206 8120 8262 8129
rect 8206 8055 8208 8064
rect 8260 8055 8262 8064
rect 8208 8026 8260 8032
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 8116 7404 8168 7410
rect 8220 7392 8248 8026
rect 8404 7546 8432 8298
rect 8588 7954 8616 8434
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8588 7478 8616 7890
rect 8576 7472 8628 7478
rect 8576 7414 8628 7420
rect 8168 7364 8248 7392
rect 8300 7404 8352 7410
rect 8116 7346 8168 7352
rect 8300 7346 8352 7352
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7760 5914 7788 6258
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 8116 3732 8168 3738
rect 8312 3720 8340 7346
rect 8392 6724 8444 6730
rect 8392 6666 8444 6672
rect 8404 6458 8432 6666
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8484 6384 8536 6390
rect 8484 6326 8536 6332
rect 8496 4146 8524 6326
rect 8772 5302 8800 8434
rect 8760 5296 8812 5302
rect 8760 5238 8812 5244
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8168 3692 8340 3720
rect 8116 3674 8168 3680
rect 8496 3670 8524 4082
rect 7564 3664 7616 3670
rect 7564 3606 7616 3612
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 5000 800 5028 2382
rect 5368 800 5396 2790
rect 6104 800 6132 2994
rect 6472 800 6500 3470
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 6840 800 6868 2246
rect 6932 2106 6960 2382
rect 6920 2100 6972 2106
rect 6920 2042 6972 2048
rect 7576 800 7604 2382
rect 7944 800 7972 3470
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8312 3058 8340 3334
rect 8772 3126 8800 5238
rect 8864 3942 8892 9438
rect 9140 9178 9168 9998
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 8944 9104 8996 9110
rect 8944 9046 8996 9052
rect 8956 8974 8984 9046
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 8956 7342 8984 8910
rect 9140 8634 9168 8910
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9232 8498 9260 11766
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9416 7546 9444 8230
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8956 6798 8984 7278
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 9312 6724 9364 6730
rect 9312 6666 9364 6672
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 9140 5778 9168 6394
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9324 4622 9352 6666
rect 9508 5370 9536 7686
rect 9600 6866 9628 8978
rect 9876 8838 9904 22066
rect 10612 22066 10732 22094
rect 10416 20868 10468 20874
rect 10416 20810 10468 20816
rect 10428 20602 10456 20810
rect 10416 20596 10468 20602
rect 10416 20538 10468 20544
rect 10508 18760 10560 18766
rect 10508 18702 10560 18708
rect 9956 17536 10008 17542
rect 9956 17478 10008 17484
rect 9968 9674 9996 17478
rect 10520 16046 10548 18702
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10336 15502 10364 15846
rect 10520 15502 10548 15982
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10612 14890 10640 22066
rect 10876 22024 10928 22030
rect 10876 21966 10928 21972
rect 10888 21486 10916 21966
rect 11256 21894 11284 22578
rect 11336 21956 11388 21962
rect 11336 21898 11388 21904
rect 11244 21888 11296 21894
rect 11244 21830 11296 21836
rect 10876 21480 10928 21486
rect 10876 21422 10928 21428
rect 10888 19854 10916 21422
rect 11348 21146 11376 21898
rect 11336 21140 11388 21146
rect 11336 21082 11388 21088
rect 10876 19848 10928 19854
rect 10876 19790 10928 19796
rect 10888 19514 10916 19790
rect 11060 19780 11112 19786
rect 11060 19722 11112 19728
rect 10876 19508 10928 19514
rect 10876 19450 10928 19456
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 10796 18426 10824 19314
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10692 16720 10744 16726
rect 10692 16662 10744 16668
rect 10704 15978 10732 16662
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10692 15972 10744 15978
rect 10692 15914 10744 15920
rect 10796 15638 10824 16050
rect 10888 15706 10916 19450
rect 11072 18970 11100 19722
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 11060 18964 11112 18970
rect 11060 18906 11112 18912
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 10968 18624 11020 18630
rect 10968 18566 11020 18572
rect 10980 18154 11008 18566
rect 10968 18148 11020 18154
rect 10968 18090 11020 18096
rect 10968 17672 11020 17678
rect 11072 17660 11100 18702
rect 11164 17814 11192 19110
rect 11152 17808 11204 17814
rect 11152 17750 11204 17756
rect 11164 17678 11192 17750
rect 11020 17632 11100 17660
rect 11152 17672 11204 17678
rect 10968 17614 11020 17620
rect 11152 17614 11204 17620
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 10980 16590 11008 17614
rect 11348 16697 11376 17614
rect 11334 16688 11390 16697
rect 11334 16623 11336 16632
rect 11388 16623 11390 16632
rect 11336 16594 11388 16600
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 11244 16584 11296 16590
rect 11348 16563 11376 16594
rect 11244 16526 11296 16532
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10784 15632 10836 15638
rect 10784 15574 10836 15580
rect 10600 14884 10652 14890
rect 10600 14826 10652 14832
rect 10324 14272 10376 14278
rect 10324 14214 10376 14220
rect 10048 14000 10100 14006
rect 10048 13942 10100 13948
rect 10060 12782 10088 13942
rect 10336 13870 10364 14214
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10324 13252 10376 13258
rect 10324 13194 10376 13200
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 10244 12782 10272 13126
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 10244 12238 10272 12582
rect 10336 12442 10364 13194
rect 10428 12714 10456 13670
rect 10416 12708 10468 12714
rect 10416 12650 10468 12656
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10428 11150 10456 12174
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 10048 11008 10100 11014
rect 10048 10950 10100 10956
rect 10060 10674 10088 10950
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10336 10674 10364 10746
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 9968 9646 10364 9674
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10152 8906 10180 9318
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9692 7886 9720 8774
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 9876 7886 9904 8366
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9600 6390 9628 6802
rect 9956 6724 10008 6730
rect 9956 6666 10008 6672
rect 9588 6384 9640 6390
rect 9588 6326 9640 6332
rect 9968 5914 9996 6666
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 9588 5840 9640 5846
rect 9588 5782 9640 5788
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9128 4616 9180 4622
rect 9048 4576 9128 4604
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8956 3602 8984 3878
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 9048 3534 9076 4576
rect 9128 4558 9180 4564
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 9140 4214 9168 4422
rect 9128 4208 9180 4214
rect 9128 4150 9180 4156
rect 9600 4146 9628 5782
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9600 3738 9628 4082
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 9632 3598 9688 3607
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 9140 3194 9168 3538
rect 9632 3533 9688 3542
rect 9864 3528 9916 3534
rect 9770 3496 9826 3505
rect 9864 3470 9916 3476
rect 9770 3431 9772 3440
rect 9824 3431 9826 3440
rect 9772 3402 9824 3408
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9692 3194 9720 3334
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 9692 2774 9720 2858
rect 9876 2854 9904 3470
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 9968 3058 9996 3334
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 9416 2746 9720 2774
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 8300 2304 8352 2310
rect 8300 2246 8352 2252
rect 8312 800 8340 2246
rect 8956 2038 8984 2382
rect 9036 2372 9088 2378
rect 9036 2314 9088 2320
rect 8944 2032 8996 2038
rect 8944 1974 8996 1980
rect 9048 800 9076 2314
rect 9416 800 9444 2746
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 9784 800 9812 2246
rect 10152 800 10180 4558
rect 10244 2922 10272 5170
rect 10232 2916 10284 2922
rect 10232 2858 10284 2864
rect 10336 2446 10364 9646
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10428 6322 10456 6598
rect 10416 6316 10468 6322
rect 10416 6258 10468 6264
rect 10416 5636 10468 5642
rect 10416 5578 10468 5584
rect 10428 4826 10456 5578
rect 10520 5370 10548 13874
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10612 10198 10640 10474
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 10704 10130 10732 12718
rect 10876 12708 10928 12714
rect 10876 12650 10928 12656
rect 10888 11898 10916 12650
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10784 11076 10836 11082
rect 10784 11018 10836 11024
rect 10796 10470 10824 11018
rect 10888 10538 10916 11834
rect 10876 10532 10928 10538
rect 10876 10474 10928 10480
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10888 10062 10916 10474
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10612 5710 10640 6734
rect 10692 6384 10744 6390
rect 10692 6326 10744 6332
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10428 4010 10456 4762
rect 10416 4004 10468 4010
rect 10416 3946 10468 3952
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10520 800 10548 5170
rect 10600 4548 10652 4554
rect 10600 4490 10652 4496
rect 10612 3942 10640 4490
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10704 3505 10732 6326
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10796 5710 10824 6054
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10690 3496 10746 3505
rect 10690 3431 10746 3440
rect 10600 2848 10652 2854
rect 10600 2790 10652 2796
rect 10612 2310 10640 2790
rect 10600 2304 10652 2310
rect 10600 2246 10652 2252
rect 10876 2304 10928 2310
rect 10876 2246 10928 2252
rect 10888 800 10916 2246
rect 10980 2106 11008 16390
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 11164 15706 11192 15982
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11256 15638 11284 16526
rect 11244 15632 11296 15638
rect 11244 15574 11296 15580
rect 11440 10606 11468 23666
rect 11532 22710 11560 23802
rect 11716 23798 11744 25094
rect 12176 24886 12204 25094
rect 12164 24880 12216 24886
rect 12164 24822 12216 24828
rect 11796 24132 11848 24138
rect 11796 24074 11848 24080
rect 11704 23792 11756 23798
rect 11704 23734 11756 23740
rect 11716 23322 11744 23734
rect 11704 23316 11756 23322
rect 11704 23258 11756 23264
rect 11716 22710 11744 23258
rect 11808 23118 11836 24074
rect 11796 23112 11848 23118
rect 11796 23054 11848 23060
rect 11520 22704 11572 22710
rect 11520 22646 11572 22652
rect 11704 22704 11756 22710
rect 11704 22646 11756 22652
rect 11532 21962 11560 22646
rect 11520 21956 11572 21962
rect 11520 21898 11572 21904
rect 11520 20460 11572 20466
rect 11520 20402 11572 20408
rect 11532 17882 11560 20402
rect 11704 19780 11756 19786
rect 11704 19722 11756 19728
rect 11716 19310 11744 19722
rect 11704 19304 11756 19310
rect 11704 19246 11756 19252
rect 11716 18290 11744 19246
rect 11612 18284 11664 18290
rect 11612 18226 11664 18232
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 11624 17882 11652 18226
rect 11520 17876 11572 17882
rect 11520 17818 11572 17824
rect 11612 17876 11664 17882
rect 11612 17818 11664 17824
rect 11612 15428 11664 15434
rect 11716 15416 11744 18226
rect 11808 16250 11836 23054
rect 12360 22982 12388 28966
rect 12532 25832 12584 25838
rect 12532 25774 12584 25780
rect 12348 22976 12400 22982
rect 12348 22918 12400 22924
rect 12440 22568 12492 22574
rect 12440 22510 12492 22516
rect 12164 22500 12216 22506
rect 12164 22442 12216 22448
rect 11888 22432 11940 22438
rect 11888 22374 11940 22380
rect 11900 20942 11928 22374
rect 12176 22234 12204 22442
rect 12348 22432 12400 22438
rect 12348 22374 12400 22380
rect 12164 22228 12216 22234
rect 12164 22170 12216 22176
rect 12360 21622 12388 22374
rect 12452 22030 12480 22510
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12348 21616 12400 21622
rect 12348 21558 12400 21564
rect 11888 20936 11940 20942
rect 11888 20878 11940 20884
rect 12348 19712 12400 19718
rect 12348 19654 12400 19660
rect 12072 18760 12124 18766
rect 12072 18702 12124 18708
rect 11980 18692 12032 18698
rect 11980 18634 12032 18640
rect 11992 18426 12020 18634
rect 11980 18420 12032 18426
rect 11980 18362 12032 18368
rect 11980 17672 12032 17678
rect 12084 17660 12112 18702
rect 12256 18624 12308 18630
rect 12256 18566 12308 18572
rect 12032 17632 12112 17660
rect 11980 17614 12032 17620
rect 12072 17536 12124 17542
rect 12072 17478 12124 17484
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 11664 15388 11744 15416
rect 11612 15370 11664 15376
rect 11624 15094 11652 15370
rect 11612 15088 11664 15094
rect 11612 15030 11664 15036
rect 11808 15026 11836 16186
rect 12084 15502 12112 17478
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 11612 14340 11664 14346
rect 11612 14282 11664 14288
rect 11624 14074 11652 14282
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11808 12782 11836 13874
rect 12084 13394 12112 14350
rect 12164 14000 12216 14006
rect 12164 13942 12216 13948
rect 12176 13802 12204 13942
rect 12164 13796 12216 13802
rect 12164 13738 12216 13744
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11808 12238 11836 12718
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 12176 12170 12204 13738
rect 12164 12164 12216 12170
rect 12164 12106 12216 12112
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11532 10674 11560 11086
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11336 10056 11388 10062
rect 11256 10016 11336 10044
rect 11256 9926 11284 10016
rect 11336 9998 11388 10004
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11072 8090 11100 9522
rect 11532 9042 11560 10610
rect 11624 10266 11652 10610
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11532 8634 11560 8978
rect 11808 8974 11836 9318
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11808 8378 11836 8434
rect 11716 8350 11836 8378
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 11072 3398 11100 7278
rect 11150 6760 11206 6769
rect 11150 6695 11152 6704
rect 11204 6695 11206 6704
rect 11152 6666 11204 6672
rect 11612 6248 11664 6254
rect 11612 6190 11664 6196
rect 11624 5710 11652 6190
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 11164 3738 11192 4014
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 11164 3058 11192 3674
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 10968 2100 11020 2106
rect 10968 2042 11020 2048
rect 11256 800 11284 4558
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11348 4146 11376 4422
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11440 2514 11468 5510
rect 11716 5370 11744 8350
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11808 7886 11836 8230
rect 11992 8090 12020 9522
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 12084 7274 12112 8366
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12176 8022 12204 8230
rect 12164 8016 12216 8022
rect 12164 7958 12216 7964
rect 12072 7268 12124 7274
rect 12072 7210 12124 7216
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11808 5692 11836 6258
rect 11888 5704 11940 5710
rect 11808 5664 11888 5692
rect 11888 5646 11940 5652
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11612 5228 11664 5234
rect 11612 5170 11664 5176
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 11532 3641 11560 4150
rect 11518 3632 11574 3641
rect 11518 3567 11574 3576
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 11532 2106 11560 2382
rect 11520 2100 11572 2106
rect 11520 2042 11572 2048
rect 11624 800 11652 5170
rect 11796 4752 11848 4758
rect 11796 4694 11848 4700
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11716 3126 11744 4014
rect 11808 3126 11836 4694
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 11796 3120 11848 3126
rect 11796 3062 11848 3068
rect 11900 3058 11928 5646
rect 11992 5574 12020 6734
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 12084 3466 12112 4422
rect 12072 3460 12124 3466
rect 12072 3402 12124 3408
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 12268 2774 12296 18566
rect 12360 18358 12388 19654
rect 12348 18352 12400 18358
rect 12348 18294 12400 18300
rect 12544 17338 12572 25774
rect 12636 18834 12664 33798
rect 12716 33448 12768 33454
rect 12716 33390 12768 33396
rect 12728 32910 12756 33390
rect 12716 32904 12768 32910
rect 12716 32846 12768 32852
rect 12820 32842 12848 36654
rect 13004 35834 13032 41006
rect 13084 40928 13136 40934
rect 13084 40870 13136 40876
rect 13096 40730 13124 40870
rect 13084 40724 13136 40730
rect 13084 40666 13136 40672
rect 13188 40458 13216 41142
rect 13268 41132 13320 41138
rect 13268 41074 13320 41080
rect 13280 40934 13308 41074
rect 13268 40928 13320 40934
rect 13268 40870 13320 40876
rect 13176 40452 13228 40458
rect 13176 40394 13228 40400
rect 13084 40384 13136 40390
rect 13084 40326 13136 40332
rect 13096 39642 13124 40326
rect 13084 39636 13136 39642
rect 13084 39578 13136 39584
rect 13188 36378 13216 40394
rect 13268 40384 13320 40390
rect 13268 40326 13320 40332
rect 13280 40118 13308 40326
rect 13268 40112 13320 40118
rect 13268 40054 13320 40060
rect 13268 37256 13320 37262
rect 13268 37198 13320 37204
rect 13176 36372 13228 36378
rect 13176 36314 13228 36320
rect 13084 36168 13136 36174
rect 13084 36110 13136 36116
rect 12992 35828 13044 35834
rect 12992 35770 13044 35776
rect 12900 35760 12952 35766
rect 12900 35702 12952 35708
rect 12912 35086 12940 35702
rect 12992 35624 13044 35630
rect 12992 35566 13044 35572
rect 13004 35193 13032 35566
rect 12990 35184 13046 35193
rect 12990 35119 13046 35128
rect 12900 35080 12952 35086
rect 12900 35022 12952 35028
rect 12992 35012 13044 35018
rect 12992 34954 13044 34960
rect 12900 34672 12952 34678
rect 12900 34614 12952 34620
rect 12808 32836 12860 32842
rect 12808 32778 12860 32784
rect 12820 31482 12848 32778
rect 12808 31476 12860 31482
rect 12808 31418 12860 31424
rect 12820 30802 12848 31418
rect 12808 30796 12860 30802
rect 12808 30738 12860 30744
rect 12714 29200 12770 29209
rect 12714 29135 12770 29144
rect 12808 29164 12860 29170
rect 12728 28490 12756 29135
rect 12808 29106 12860 29112
rect 12820 28762 12848 29106
rect 12808 28756 12860 28762
rect 12808 28698 12860 28704
rect 12716 28484 12768 28490
rect 12716 28426 12768 28432
rect 12716 27940 12768 27946
rect 12716 27882 12768 27888
rect 12728 27470 12756 27882
rect 12716 27464 12768 27470
rect 12716 27406 12768 27412
rect 12912 26586 12940 34614
rect 13004 30054 13032 34954
rect 13096 33930 13124 36110
rect 13176 35080 13228 35086
rect 13176 35022 13228 35028
rect 13084 33924 13136 33930
rect 13084 33866 13136 33872
rect 12992 30048 13044 30054
rect 12992 29990 13044 29996
rect 13096 29714 13124 33866
rect 13084 29708 13136 29714
rect 13084 29650 13136 29656
rect 13188 29594 13216 35022
rect 13280 33046 13308 37198
rect 13372 33998 13400 41386
rect 13450 41304 13506 41313
rect 13450 41239 13506 41248
rect 13464 41002 13492 41239
rect 13452 40996 13504 41002
rect 13452 40938 13504 40944
rect 13452 38208 13504 38214
rect 13452 38150 13504 38156
rect 13464 37466 13492 38150
rect 13452 37460 13504 37466
rect 13452 37402 13504 37408
rect 13556 37126 13584 45358
rect 13924 45354 13952 45834
rect 14016 45490 14044 46514
rect 14476 46170 14504 46514
rect 14844 46442 14872 46990
rect 15120 46510 15148 48010
rect 15396 47258 15424 49200
rect 15384 47252 15436 47258
rect 15384 47194 15436 47200
rect 15568 47048 15620 47054
rect 15568 46990 15620 46996
rect 15580 46714 15608 46990
rect 16224 46918 16252 49200
rect 16304 47728 16356 47734
rect 16304 47670 16356 47676
rect 16212 46912 16264 46918
rect 16212 46854 16264 46860
rect 15568 46708 15620 46714
rect 15568 46650 15620 46656
rect 15108 46504 15160 46510
rect 15108 46446 15160 46452
rect 14832 46436 14884 46442
rect 14832 46378 14884 46384
rect 14924 46368 14976 46374
rect 14924 46310 14976 46316
rect 14936 46170 14964 46310
rect 14464 46164 14516 46170
rect 14464 46106 14516 46112
rect 14924 46164 14976 46170
rect 14924 46106 14976 46112
rect 14096 46028 14148 46034
rect 14096 45970 14148 45976
rect 15108 46028 15160 46034
rect 15108 45970 15160 45976
rect 14004 45484 14056 45490
rect 14004 45426 14056 45432
rect 13912 45348 13964 45354
rect 13912 45290 13964 45296
rect 14108 43466 14136 45970
rect 14464 45960 14516 45966
rect 14464 45902 14516 45908
rect 14476 44198 14504 45902
rect 14556 44396 14608 44402
rect 14556 44338 14608 44344
rect 14832 44396 14884 44402
rect 14832 44338 14884 44344
rect 14464 44192 14516 44198
rect 14464 44134 14516 44140
rect 14476 43790 14504 44134
rect 14464 43784 14516 43790
rect 14464 43726 14516 43732
rect 14016 43450 14136 43466
rect 14016 43444 14148 43450
rect 14016 43438 14096 43444
rect 14016 42702 14044 43438
rect 14096 43386 14148 43392
rect 14096 43308 14148 43314
rect 14096 43250 14148 43256
rect 14108 42770 14136 43250
rect 14096 42764 14148 42770
rect 14096 42706 14148 42712
rect 14188 42764 14240 42770
rect 14188 42706 14240 42712
rect 14004 42696 14056 42702
rect 14004 42638 14056 42644
rect 14016 42566 14044 42638
rect 14004 42560 14056 42566
rect 14004 42502 14056 42508
rect 14200 42158 14228 42706
rect 14372 42696 14424 42702
rect 14372 42638 14424 42644
rect 14280 42220 14332 42226
rect 14280 42162 14332 42168
rect 14188 42152 14240 42158
rect 14188 42094 14240 42100
rect 14200 41682 14228 42094
rect 14188 41676 14240 41682
rect 14188 41618 14240 41624
rect 13728 41064 13780 41070
rect 13728 41006 13780 41012
rect 13740 40769 13768 41006
rect 13726 40760 13782 40769
rect 13726 40695 13782 40704
rect 14188 39840 14240 39846
rect 14188 39782 14240 39788
rect 14096 37936 14148 37942
rect 14096 37878 14148 37884
rect 13636 37868 13688 37874
rect 13636 37810 13688 37816
rect 13648 37194 13676 37810
rect 13728 37732 13780 37738
rect 13728 37674 13780 37680
rect 13740 37398 13768 37674
rect 13728 37392 13780 37398
rect 13728 37334 13780 37340
rect 13636 37188 13688 37194
rect 13636 37130 13688 37136
rect 13544 37120 13596 37126
rect 13544 37062 13596 37068
rect 13648 36938 13676 37130
rect 13556 36910 13676 36938
rect 13740 36922 13768 37334
rect 14108 36922 14136 37878
rect 13728 36916 13780 36922
rect 13360 33992 13412 33998
rect 13412 33952 13492 33980
rect 13360 33934 13412 33940
rect 13268 33040 13320 33046
rect 13268 32982 13320 32988
rect 13360 32904 13412 32910
rect 13360 32846 13412 32852
rect 13268 32428 13320 32434
rect 13268 32370 13320 32376
rect 13280 30734 13308 32370
rect 13268 30728 13320 30734
rect 13268 30670 13320 30676
rect 13372 30546 13400 32846
rect 13004 29566 13216 29594
rect 13280 30518 13400 30546
rect 12900 26580 12952 26586
rect 12900 26522 12952 26528
rect 12808 25696 12860 25702
rect 12808 25638 12860 25644
rect 12820 25294 12848 25638
rect 12900 25492 12952 25498
rect 12900 25434 12952 25440
rect 12808 25288 12860 25294
rect 12808 25230 12860 25236
rect 12820 24274 12848 25230
rect 12912 24954 12940 25434
rect 12900 24948 12952 24954
rect 12900 24890 12952 24896
rect 12808 24268 12860 24274
rect 12728 24228 12808 24256
rect 12728 21146 12756 24228
rect 12808 24210 12860 24216
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 12912 22234 12940 22578
rect 12808 22228 12860 22234
rect 12808 22170 12860 22176
rect 12900 22228 12952 22234
rect 12900 22170 12952 22176
rect 12820 21690 12848 22170
rect 12900 22094 12952 22098
rect 13004 22094 13032 29566
rect 13176 29504 13228 29510
rect 13176 29446 13228 29452
rect 13084 29300 13136 29306
rect 13084 29242 13136 29248
rect 13096 25650 13124 29242
rect 13188 28558 13216 29446
rect 13176 28552 13228 28558
rect 13176 28494 13228 28500
rect 13176 27396 13228 27402
rect 13176 27338 13228 27344
rect 13188 27169 13216 27338
rect 13174 27160 13230 27169
rect 13174 27095 13230 27104
rect 13176 26920 13228 26926
rect 13176 26862 13228 26868
rect 13188 25838 13216 26862
rect 13280 26518 13308 30518
rect 13464 30394 13492 33952
rect 13556 33590 13584 36910
rect 13728 36858 13780 36864
rect 14096 36916 14148 36922
rect 14096 36858 14148 36864
rect 13820 36712 13872 36718
rect 13820 36654 13872 36660
rect 13728 34740 13780 34746
rect 13728 34682 13780 34688
rect 13636 34604 13688 34610
rect 13636 34546 13688 34552
rect 13648 33658 13676 34546
rect 13636 33652 13688 33658
rect 13636 33594 13688 33600
rect 13544 33584 13596 33590
rect 13544 33526 13596 33532
rect 13634 33552 13690 33561
rect 13634 33487 13636 33496
rect 13688 33487 13690 33496
rect 13636 33458 13688 33464
rect 13648 32978 13676 33458
rect 13636 32972 13688 32978
rect 13636 32914 13688 32920
rect 13636 32224 13688 32230
rect 13636 32166 13688 32172
rect 13648 31890 13676 32166
rect 13636 31884 13688 31890
rect 13636 31826 13688 31832
rect 13636 31680 13688 31686
rect 13636 31622 13688 31628
rect 13648 31482 13676 31622
rect 13636 31476 13688 31482
rect 13636 31418 13688 31424
rect 13544 31340 13596 31346
rect 13544 31282 13596 31288
rect 13556 30938 13584 31282
rect 13648 30938 13676 31418
rect 13544 30932 13596 30938
rect 13544 30874 13596 30880
rect 13636 30932 13688 30938
rect 13636 30874 13688 30880
rect 13544 30796 13596 30802
rect 13544 30738 13596 30744
rect 13636 30796 13688 30802
rect 13636 30738 13688 30744
rect 13452 30388 13504 30394
rect 13452 30330 13504 30336
rect 13556 30274 13584 30738
rect 13648 30326 13676 30738
rect 13372 30246 13584 30274
rect 13636 30320 13688 30326
rect 13636 30262 13688 30268
rect 13268 26512 13320 26518
rect 13268 26454 13320 26460
rect 13268 26376 13320 26382
rect 13268 26318 13320 26324
rect 13280 26042 13308 26318
rect 13268 26036 13320 26042
rect 13268 25978 13320 25984
rect 13372 25838 13400 30246
rect 13636 30048 13688 30054
rect 13636 29990 13688 29996
rect 13452 29708 13504 29714
rect 13452 29650 13504 29656
rect 13176 25832 13228 25838
rect 13360 25832 13412 25838
rect 13176 25774 13228 25780
rect 13358 25800 13360 25809
rect 13412 25800 13414 25809
rect 13358 25735 13414 25744
rect 13096 25622 13308 25650
rect 13280 23594 13308 25622
rect 13360 24744 13412 24750
rect 13360 24686 13412 24692
rect 13372 23733 13400 24686
rect 13357 23727 13409 23733
rect 13357 23669 13409 23675
rect 13268 23588 13320 23594
rect 13268 23530 13320 23536
rect 13084 23520 13136 23526
rect 13084 23462 13136 23468
rect 13096 22642 13124 23462
rect 13084 22636 13136 22642
rect 13084 22578 13136 22584
rect 13084 22228 13136 22234
rect 13084 22170 13136 22176
rect 12900 22092 13032 22094
rect 12952 22066 13032 22092
rect 12900 22034 12952 22040
rect 12808 21684 12860 21690
rect 12808 21626 12860 21632
rect 12716 21140 12768 21146
rect 12716 21082 12768 21088
rect 12728 19334 12756 21082
rect 12912 20942 12940 22034
rect 13096 21894 13124 22170
rect 13084 21888 13136 21894
rect 13084 21830 13136 21836
rect 12900 20936 12952 20942
rect 12900 20878 12952 20884
rect 12912 20602 12940 20878
rect 12900 20596 12952 20602
rect 12900 20538 12952 20544
rect 12728 19306 12848 19334
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 12820 17746 12848 19306
rect 13176 18760 13228 18766
rect 13176 18702 13228 18708
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 12912 18057 12940 18566
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 12898 18048 12954 18057
rect 12898 17983 12954 17992
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 12624 17672 12676 17678
rect 12624 17614 12676 17620
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12452 13870 12480 14554
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12544 12434 12572 17274
rect 12636 17066 12664 17614
rect 13096 17542 13124 18226
rect 13188 17882 13216 18702
rect 13280 17954 13308 23530
rect 13464 23050 13492 29650
rect 13544 29640 13596 29646
rect 13544 29582 13596 29588
rect 13556 28218 13584 29582
rect 13648 29578 13676 29990
rect 13636 29572 13688 29578
rect 13636 29514 13688 29520
rect 13544 28212 13596 28218
rect 13544 28154 13596 28160
rect 13544 27328 13596 27334
rect 13544 27270 13596 27276
rect 13556 24886 13584 27270
rect 13544 24880 13596 24886
rect 13544 24822 13596 24828
rect 13648 24818 13676 29514
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13452 23044 13504 23050
rect 13452 22986 13504 22992
rect 13464 22778 13492 22986
rect 13452 22772 13504 22778
rect 13452 22714 13504 22720
rect 13280 17926 13400 17954
rect 13176 17876 13228 17882
rect 13176 17818 13228 17824
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 12992 17332 13044 17338
rect 12992 17274 13044 17280
rect 12624 17060 12676 17066
rect 12624 17002 12676 17008
rect 12636 16182 12664 17002
rect 12624 16176 12676 16182
rect 12624 16118 12676 16124
rect 12636 15586 12664 16118
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12728 15706 12756 16050
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12636 15558 12756 15586
rect 12728 15434 12756 15558
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 12716 15428 12768 15434
rect 12716 15370 12768 15376
rect 12728 12434 12756 15370
rect 12912 15366 12940 15438
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 12912 12918 12940 13194
rect 12900 12912 12952 12918
rect 12900 12854 12952 12860
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12820 12753 12848 12786
rect 12806 12744 12862 12753
rect 12806 12679 12862 12688
rect 13004 12434 13032 17274
rect 13096 17270 13124 17478
rect 13084 17264 13136 17270
rect 13084 17206 13136 17212
rect 13084 16584 13136 16590
rect 13188 16572 13216 17818
rect 13136 16544 13216 16572
rect 13268 16562 13320 16568
rect 13084 16526 13136 16532
rect 13268 16504 13320 16510
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 12452 12406 12572 12434
rect 12636 12406 12756 12434
rect 12820 12406 13032 12434
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12360 11150 12388 11494
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12452 9654 12480 12406
rect 12636 11762 12664 12406
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12636 9586 12664 11698
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12728 10062 12756 11494
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12360 7954 12388 8910
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 12728 7410 12756 9454
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12544 6390 12572 6598
rect 12532 6384 12584 6390
rect 12532 6326 12584 6332
rect 12820 6254 12848 12406
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 12912 10538 12940 11630
rect 12900 10532 12952 10538
rect 12900 10474 12952 10480
rect 12912 10130 12940 10474
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 13004 8498 13032 9318
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 12992 8016 13044 8022
rect 12992 7958 13044 7964
rect 13004 7478 13032 7958
rect 12992 7472 13044 7478
rect 12992 7414 13044 7420
rect 12992 6860 13044 6866
rect 12992 6802 13044 6808
rect 12898 6760 12954 6769
rect 12898 6695 12900 6704
rect 12952 6695 12954 6704
rect 12900 6666 12952 6672
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12452 5166 12480 6054
rect 12728 5846 12756 6054
rect 12716 5840 12768 5846
rect 12716 5782 12768 5788
rect 12820 5710 12848 6190
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12452 3194 12480 4558
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12544 3738 12572 4082
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12360 2990 12388 3130
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12636 2854 12664 4558
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12820 4214 12848 4422
rect 12808 4208 12860 4214
rect 12808 4150 12860 4156
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12728 3058 12756 3878
rect 12716 3052 12768 3058
rect 12716 2994 12768 3000
rect 12348 2848 12400 2854
rect 12348 2790 12400 2796
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 12176 2746 12296 2774
rect 12176 2582 12204 2746
rect 12164 2576 12216 2582
rect 12164 2518 12216 2524
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 11992 800 12020 2246
rect 12360 800 12388 2790
rect 12912 2774 12940 6258
rect 13004 5778 13032 6802
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 13004 3602 13032 5714
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 13004 3126 13032 3538
rect 12992 3120 13044 3126
rect 12992 3062 13044 3068
rect 13096 2774 13124 16390
rect 13188 15502 13216 16390
rect 13280 15570 13308 16504
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 13176 15496 13228 15502
rect 13176 15438 13228 15444
rect 13188 15144 13216 15438
rect 13268 15156 13320 15162
rect 13188 15116 13268 15144
rect 13268 15098 13320 15104
rect 13176 14340 13228 14346
rect 13176 14282 13228 14288
rect 13188 14074 13216 14282
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 13176 13796 13228 13802
rect 13176 13738 13228 13744
rect 13188 6458 13216 13738
rect 13280 12850 13308 13874
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 13372 9382 13400 17926
rect 13452 17740 13504 17746
rect 13452 17682 13504 17688
rect 13464 17338 13492 17682
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13464 15978 13492 16390
rect 13452 15972 13504 15978
rect 13452 15914 13504 15920
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13556 15094 13584 15846
rect 13544 15088 13596 15094
rect 13544 15030 13596 15036
rect 13648 13530 13676 24754
rect 13740 16794 13768 34682
rect 13832 33862 13860 36654
rect 14004 35488 14056 35494
rect 14004 35430 14056 35436
rect 13912 34740 13964 34746
rect 13912 34682 13964 34688
rect 13820 33856 13872 33862
rect 13820 33798 13872 33804
rect 13832 32366 13860 33798
rect 13820 32360 13872 32366
rect 13820 32302 13872 32308
rect 13832 32026 13860 32302
rect 13820 32020 13872 32026
rect 13820 31962 13872 31968
rect 13820 31476 13872 31482
rect 13820 31418 13872 31424
rect 13832 31346 13860 31418
rect 13820 31340 13872 31346
rect 13820 31282 13872 31288
rect 13820 30320 13872 30326
rect 13820 30262 13872 30268
rect 13832 27334 13860 30262
rect 13820 27328 13872 27334
rect 13820 27270 13872 27276
rect 13820 26920 13872 26926
rect 13820 26862 13872 26868
rect 13832 25906 13860 26862
rect 13820 25900 13872 25906
rect 13820 25842 13872 25848
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 13832 24342 13860 24754
rect 13820 24336 13872 24342
rect 13820 24278 13872 24284
rect 13924 24154 13952 34682
rect 14016 25838 14044 35430
rect 14096 35284 14148 35290
rect 14096 35226 14148 35232
rect 14108 29306 14136 35226
rect 14200 35086 14228 39782
rect 14292 39370 14320 42162
rect 14384 42022 14412 42638
rect 14372 42016 14424 42022
rect 14372 41958 14424 41964
rect 14280 39364 14332 39370
rect 14280 39306 14332 39312
rect 14280 38344 14332 38350
rect 14280 38286 14332 38292
rect 14292 38010 14320 38286
rect 14372 38208 14424 38214
rect 14372 38150 14424 38156
rect 14280 38004 14332 38010
rect 14280 37946 14332 37952
rect 14384 37194 14412 38150
rect 14372 37188 14424 37194
rect 14372 37130 14424 37136
rect 14280 35828 14332 35834
rect 14280 35770 14332 35776
rect 14188 35080 14240 35086
rect 14188 35022 14240 35028
rect 14292 34542 14320 35770
rect 14476 35222 14504 43726
rect 14568 43450 14596 44338
rect 14648 44328 14700 44334
rect 14648 44270 14700 44276
rect 14660 43790 14688 44270
rect 14648 43784 14700 43790
rect 14648 43726 14700 43732
rect 14556 43444 14608 43450
rect 14556 43386 14608 43392
rect 14660 43382 14688 43726
rect 14648 43376 14700 43382
rect 14648 43318 14700 43324
rect 14556 41540 14608 41546
rect 14556 41482 14608 41488
rect 14464 35216 14516 35222
rect 14464 35158 14516 35164
rect 14568 35034 14596 41482
rect 14660 40594 14688 43318
rect 14740 42696 14792 42702
rect 14740 42638 14792 42644
rect 14752 42242 14780 42638
rect 14844 42362 14872 44338
rect 15016 43648 15068 43654
rect 15016 43590 15068 43596
rect 15028 43314 15056 43590
rect 14924 43308 14976 43314
rect 14924 43250 14976 43256
rect 15016 43308 15068 43314
rect 15016 43250 15068 43256
rect 14936 42770 14964 43250
rect 14924 42764 14976 42770
rect 14924 42706 14976 42712
rect 14924 42560 14976 42566
rect 14924 42502 14976 42508
rect 14832 42356 14884 42362
rect 14832 42298 14884 42304
rect 14752 42226 14872 42242
rect 14752 42220 14884 42226
rect 14752 42214 14832 42220
rect 14832 42162 14884 42168
rect 14844 42022 14872 42162
rect 14740 42016 14792 42022
rect 14740 41958 14792 41964
rect 14832 42016 14884 42022
rect 14832 41958 14884 41964
rect 14648 40588 14700 40594
rect 14648 40530 14700 40536
rect 14648 38276 14700 38282
rect 14648 38218 14700 38224
rect 14660 37942 14688 38218
rect 14648 37936 14700 37942
rect 14648 37878 14700 37884
rect 14660 37194 14688 37878
rect 14648 37188 14700 37194
rect 14648 37130 14700 37136
rect 14372 35012 14424 35018
rect 14372 34954 14424 34960
rect 14476 35006 14596 35034
rect 14648 35080 14700 35086
rect 14648 35022 14700 35028
rect 14280 34536 14332 34542
rect 14280 34478 14332 34484
rect 14292 33980 14320 34478
rect 14384 34474 14412 34954
rect 14372 34468 14424 34474
rect 14372 34410 14424 34416
rect 14384 34082 14412 34410
rect 14476 34202 14504 35006
rect 14556 34944 14608 34950
rect 14556 34886 14608 34892
rect 14464 34196 14516 34202
rect 14464 34138 14516 34144
rect 14384 34066 14504 34082
rect 14384 34060 14516 34066
rect 14384 34054 14464 34060
rect 14464 34002 14516 34008
rect 14292 33952 14412 33980
rect 14280 33856 14332 33862
rect 14280 33798 14332 33804
rect 14292 33590 14320 33798
rect 14280 33584 14332 33590
rect 14280 33526 14332 33532
rect 14280 33312 14332 33318
rect 14278 33280 14280 33289
rect 14332 33280 14334 33289
rect 14278 33215 14334 33224
rect 14188 32904 14240 32910
rect 14188 32846 14240 32852
rect 14200 32026 14228 32846
rect 14188 32020 14240 32026
rect 14188 31962 14240 31968
rect 14200 31346 14228 31962
rect 14384 31754 14412 33952
rect 14476 32502 14504 34002
rect 14464 32496 14516 32502
rect 14464 32438 14516 32444
rect 14384 31726 14504 31754
rect 14188 31340 14240 31346
rect 14188 31282 14240 31288
rect 14372 31340 14424 31346
rect 14372 31282 14424 31288
rect 14384 30938 14412 31282
rect 14372 30932 14424 30938
rect 14372 30874 14424 30880
rect 14280 30660 14332 30666
rect 14280 30602 14332 30608
rect 14292 29646 14320 30602
rect 14280 29640 14332 29646
rect 14280 29582 14332 29588
rect 14096 29300 14148 29306
rect 14096 29242 14148 29248
rect 14108 28626 14136 29242
rect 14188 28960 14240 28966
rect 14186 28928 14188 28937
rect 14240 28928 14242 28937
rect 14186 28863 14242 28872
rect 14096 28620 14148 28626
rect 14096 28562 14148 28568
rect 14200 28558 14228 28863
rect 14188 28552 14240 28558
rect 14188 28494 14240 28500
rect 14372 27872 14424 27878
rect 14372 27814 14424 27820
rect 14280 27600 14332 27606
rect 14280 27542 14332 27548
rect 14096 27464 14148 27470
rect 14096 27406 14148 27412
rect 14108 26382 14136 27406
rect 14292 27130 14320 27542
rect 14384 27402 14412 27814
rect 14372 27396 14424 27402
rect 14372 27338 14424 27344
rect 14280 27124 14332 27130
rect 14280 27066 14332 27072
rect 14372 26988 14424 26994
rect 14372 26930 14424 26936
rect 14280 26784 14332 26790
rect 14280 26726 14332 26732
rect 14096 26376 14148 26382
rect 14096 26318 14148 26324
rect 14004 25832 14056 25838
rect 14004 25774 14056 25780
rect 14108 24614 14136 26318
rect 14188 26308 14240 26314
rect 14188 26250 14240 26256
rect 14200 26042 14228 26250
rect 14188 26036 14240 26042
rect 14188 25978 14240 25984
rect 14292 25906 14320 26726
rect 14280 25900 14332 25906
rect 14280 25842 14332 25848
rect 14188 25832 14240 25838
rect 14188 25774 14240 25780
rect 14004 24608 14056 24614
rect 14004 24550 14056 24556
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 13832 24126 13952 24154
rect 13832 20942 13860 24126
rect 14016 23798 14044 24550
rect 14004 23792 14056 23798
rect 14004 23734 14056 23740
rect 14108 23730 14136 24550
rect 13912 23724 13964 23730
rect 13912 23666 13964 23672
rect 14096 23724 14148 23730
rect 14096 23666 14148 23672
rect 13924 23633 13952 23666
rect 14004 23656 14056 23662
rect 13910 23624 13966 23633
rect 14004 23598 14056 23604
rect 13910 23559 13966 23568
rect 14016 23322 14044 23598
rect 14004 23316 14056 23322
rect 14004 23258 14056 23264
rect 14108 22030 14136 23666
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 14108 21010 14136 21966
rect 14096 21004 14148 21010
rect 14096 20946 14148 20952
rect 13820 20936 13872 20942
rect 13820 20878 13872 20884
rect 14096 20868 14148 20874
rect 14096 20810 14148 20816
rect 13820 20800 13872 20806
rect 13820 20742 13872 20748
rect 13832 20466 13860 20742
rect 13912 20596 13964 20602
rect 13912 20538 13964 20544
rect 13820 20460 13872 20466
rect 13820 20402 13872 20408
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13832 18834 13860 19654
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13832 17202 13860 17614
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13464 11286 13492 11494
rect 13452 11280 13504 11286
rect 13452 11222 13504 11228
rect 13556 9586 13584 11698
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 13832 10470 13860 11018
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13832 10062 13860 10406
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13280 8906 13308 9318
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13280 2990 13308 8842
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13372 6798 13400 7142
rect 13464 6866 13492 7346
rect 13556 7342 13584 8502
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13556 5166 13584 7278
rect 13832 6390 13860 9998
rect 13924 9110 13952 20538
rect 14004 19780 14056 19786
rect 14004 19722 14056 19728
rect 14016 18834 14044 19722
rect 14004 18828 14056 18834
rect 14004 18770 14056 18776
rect 14004 18692 14056 18698
rect 14004 18634 14056 18640
rect 14016 16590 14044 18634
rect 14004 16584 14056 16590
rect 14004 16526 14056 16532
rect 14108 15570 14136 20810
rect 14200 17218 14228 25774
rect 14280 24812 14332 24818
rect 14280 24754 14332 24760
rect 14292 23633 14320 24754
rect 14278 23624 14334 23633
rect 14278 23559 14334 23568
rect 14384 20602 14412 26930
rect 14476 26586 14504 31726
rect 14464 26580 14516 26586
rect 14464 26522 14516 26528
rect 14476 26042 14504 26522
rect 14464 26036 14516 26042
rect 14464 25978 14516 25984
rect 14464 24744 14516 24750
rect 14464 24686 14516 24692
rect 14476 24274 14504 24686
rect 14464 24268 14516 24274
rect 14464 24210 14516 24216
rect 14372 20596 14424 20602
rect 14372 20538 14424 20544
rect 14568 19990 14596 34886
rect 14660 34610 14688 35022
rect 14648 34604 14700 34610
rect 14648 34546 14700 34552
rect 14648 33312 14700 33318
rect 14648 33254 14700 33260
rect 14660 32434 14688 33254
rect 14648 32428 14700 32434
rect 14648 32370 14700 32376
rect 14752 31890 14780 41958
rect 14844 41070 14872 41958
rect 14832 41064 14884 41070
rect 14832 41006 14884 41012
rect 14936 40610 14964 42502
rect 15120 41414 15148 45970
rect 16316 45966 16344 47670
rect 17052 47258 17080 49200
rect 17500 47796 17552 47802
rect 17500 47738 17552 47744
rect 17132 47524 17184 47530
rect 17132 47466 17184 47472
rect 17040 47252 17092 47258
rect 17040 47194 17092 47200
rect 16580 47048 16632 47054
rect 16580 46990 16632 46996
rect 16488 46572 16540 46578
rect 16488 46514 16540 46520
rect 16500 46170 16528 46514
rect 16592 46442 16620 46990
rect 16580 46436 16632 46442
rect 16580 46378 16632 46384
rect 16488 46164 16540 46170
rect 16488 46106 16540 46112
rect 17144 45966 17172 47466
rect 17408 47048 17460 47054
rect 17408 46990 17460 46996
rect 17420 46714 17448 46990
rect 17408 46708 17460 46714
rect 17408 46650 17460 46656
rect 15476 45960 15528 45966
rect 15476 45902 15528 45908
rect 16304 45960 16356 45966
rect 16304 45902 16356 45908
rect 17132 45960 17184 45966
rect 17132 45902 17184 45908
rect 15488 45830 15516 45902
rect 15476 45824 15528 45830
rect 15476 45766 15528 45772
rect 15488 45286 15516 45766
rect 15476 45280 15528 45286
rect 15476 45222 15528 45228
rect 16856 44532 16908 44538
rect 16856 44474 16908 44480
rect 16672 43784 16724 43790
rect 16672 43726 16724 43732
rect 15292 43716 15344 43722
rect 15292 43658 15344 43664
rect 15200 43308 15252 43314
rect 15200 43250 15252 43256
rect 15212 42702 15240 43250
rect 15200 42696 15252 42702
rect 15200 42638 15252 42644
rect 15304 42362 15332 43658
rect 15384 43648 15436 43654
rect 15384 43590 15436 43596
rect 15396 43314 15424 43590
rect 16684 43314 16712 43726
rect 15384 43308 15436 43314
rect 15384 43250 15436 43256
rect 16672 43308 16724 43314
rect 16672 43250 16724 43256
rect 16764 43308 16816 43314
rect 16764 43250 16816 43256
rect 15292 42356 15344 42362
rect 15292 42298 15344 42304
rect 15292 41676 15344 41682
rect 15292 41618 15344 41624
rect 15200 41540 15252 41546
rect 15200 41482 15252 41488
rect 14844 40582 14964 40610
rect 15028 41386 15148 41414
rect 14844 33590 14872 40582
rect 14924 40452 14976 40458
rect 14924 40394 14976 40400
rect 14936 39642 14964 40394
rect 14924 39636 14976 39642
rect 14924 39578 14976 39584
rect 14924 38344 14976 38350
rect 14924 38286 14976 38292
rect 14936 35018 14964 38286
rect 14924 35012 14976 35018
rect 14924 34954 14976 34960
rect 14832 33584 14884 33590
rect 14832 33526 14884 33532
rect 14922 33552 14978 33561
rect 14922 33487 14924 33496
rect 14976 33487 14978 33496
rect 14924 33458 14976 33464
rect 14832 33448 14884 33454
rect 14832 33390 14884 33396
rect 14844 33318 14872 33390
rect 15028 33386 15056 41386
rect 15108 39976 15160 39982
rect 15108 39918 15160 39924
rect 15120 35834 15148 39918
rect 15212 38418 15240 41482
rect 15304 41274 15332 41618
rect 15292 41268 15344 41274
rect 15292 41210 15344 41216
rect 15396 41206 15424 43250
rect 15936 43172 15988 43178
rect 15936 43114 15988 43120
rect 15568 42220 15620 42226
rect 15844 42220 15896 42226
rect 15620 42180 15700 42208
rect 15568 42162 15620 42168
rect 15568 41268 15620 41274
rect 15568 41210 15620 41216
rect 15384 41200 15436 41206
rect 15384 41142 15436 41148
rect 15396 40905 15424 41142
rect 15580 41041 15608 41210
rect 15566 41032 15622 41041
rect 15566 40967 15622 40976
rect 15382 40896 15438 40905
rect 15382 40831 15438 40840
rect 15672 39914 15700 42180
rect 15844 42162 15896 42168
rect 15856 41682 15884 42162
rect 15844 41676 15896 41682
rect 15844 41618 15896 41624
rect 15948 41414 15976 43114
rect 16028 43104 16080 43110
rect 16028 43046 16080 43052
rect 16040 42702 16068 43046
rect 16028 42696 16080 42702
rect 16028 42638 16080 42644
rect 16212 42696 16264 42702
rect 16212 42638 16264 42644
rect 16224 42378 16252 42638
rect 16132 42350 16252 42378
rect 16132 42226 16160 42350
rect 16304 42288 16356 42294
rect 16304 42230 16356 42236
rect 16120 42220 16172 42226
rect 16120 42162 16172 42168
rect 16212 42152 16264 42158
rect 16212 42094 16264 42100
rect 15948 41386 16068 41414
rect 15844 41200 15896 41206
rect 15842 41168 15844 41177
rect 15896 41168 15898 41177
rect 15842 41103 15898 41112
rect 15856 40934 15884 41103
rect 15934 41032 15990 41041
rect 15934 40967 15990 40976
rect 15948 40934 15976 40967
rect 15844 40928 15896 40934
rect 15844 40870 15896 40876
rect 15936 40928 15988 40934
rect 15936 40870 15988 40876
rect 15936 40520 15988 40526
rect 15936 40462 15988 40468
rect 15660 39908 15712 39914
rect 15660 39850 15712 39856
rect 15384 39840 15436 39846
rect 15384 39782 15436 39788
rect 15396 39438 15424 39782
rect 15948 39506 15976 40462
rect 15660 39500 15712 39506
rect 15660 39442 15712 39448
rect 15936 39500 15988 39506
rect 15936 39442 15988 39448
rect 15384 39432 15436 39438
rect 15384 39374 15436 39380
rect 15476 39364 15528 39370
rect 15476 39306 15528 39312
rect 15292 39296 15344 39302
rect 15292 39238 15344 39244
rect 15200 38412 15252 38418
rect 15200 38354 15252 38360
rect 15108 35828 15160 35834
rect 15108 35770 15160 35776
rect 15108 34604 15160 34610
rect 15108 34546 15160 34552
rect 15120 33862 15148 34546
rect 15108 33856 15160 33862
rect 15108 33798 15160 33804
rect 14924 33380 14976 33386
rect 14924 33322 14976 33328
rect 15016 33380 15068 33386
rect 15016 33322 15068 33328
rect 14832 33312 14884 33318
rect 14936 33289 14964 33322
rect 14832 33254 14884 33260
rect 14922 33280 14978 33289
rect 14922 33215 14978 33224
rect 14936 32910 14964 33215
rect 14924 32904 14976 32910
rect 14924 32846 14976 32852
rect 14832 32768 14884 32774
rect 14832 32710 14884 32716
rect 14844 32434 14872 32710
rect 14832 32428 14884 32434
rect 14832 32370 14884 32376
rect 15028 32366 15056 33322
rect 15120 32434 15148 33798
rect 15108 32428 15160 32434
rect 15108 32370 15160 32376
rect 15016 32360 15068 32366
rect 15016 32302 15068 32308
rect 15212 32298 15240 38354
rect 15200 32292 15252 32298
rect 15200 32234 15252 32240
rect 15200 32020 15252 32026
rect 15200 31962 15252 31968
rect 14740 31884 14792 31890
rect 14740 31826 14792 31832
rect 14648 31816 14700 31822
rect 14648 31758 14700 31764
rect 14660 31482 14688 31758
rect 14648 31476 14700 31482
rect 14648 31418 14700 31424
rect 14648 30728 14700 30734
rect 14648 30670 14700 30676
rect 14660 30326 14688 30670
rect 14648 30320 14700 30326
rect 14648 30262 14700 30268
rect 14660 29646 14688 30262
rect 14648 29640 14700 29646
rect 14648 29582 14700 29588
rect 14648 29164 14700 29170
rect 14648 29106 14700 29112
rect 14660 28762 14688 29106
rect 14648 28756 14700 28762
rect 14648 28698 14700 28704
rect 14648 27532 14700 27538
rect 14648 27474 14700 27480
rect 14660 26246 14688 27474
rect 14752 26994 14780 31826
rect 15212 30802 15240 31962
rect 15200 30796 15252 30802
rect 15120 30756 15200 30784
rect 14924 29708 14976 29714
rect 14924 29650 14976 29656
rect 14832 29504 14884 29510
rect 14832 29446 14884 29452
rect 14844 28694 14872 29446
rect 14936 28948 14964 29650
rect 15120 28994 15148 30756
rect 15200 30738 15252 30744
rect 15200 30660 15252 30666
rect 15200 30602 15252 30608
rect 15212 30326 15240 30602
rect 15200 30320 15252 30326
rect 15200 30262 15252 30268
rect 15120 28966 15240 28994
rect 15200 28960 15252 28966
rect 14936 28920 15056 28948
rect 15028 28762 15056 28920
rect 15200 28902 15252 28908
rect 15016 28756 15068 28762
rect 15016 28698 15068 28704
rect 14832 28688 14884 28694
rect 14832 28630 14884 28636
rect 14924 28076 14976 28082
rect 14924 28018 14976 28024
rect 14832 27396 14884 27402
rect 14832 27338 14884 27344
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 14648 26240 14700 26246
rect 14648 26182 14700 26188
rect 14660 25906 14688 26182
rect 14648 25900 14700 25906
rect 14648 25842 14700 25848
rect 14648 24200 14700 24206
rect 14648 24142 14700 24148
rect 14660 23798 14688 24142
rect 14648 23792 14700 23798
rect 14648 23734 14700 23740
rect 14660 23118 14688 23734
rect 14648 23112 14700 23118
rect 14648 23054 14700 23060
rect 14740 20868 14792 20874
rect 14740 20810 14792 20816
rect 14752 20602 14780 20810
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14556 19984 14608 19990
rect 14556 19926 14608 19932
rect 14280 19780 14332 19786
rect 14280 19722 14332 19728
rect 14292 19514 14320 19722
rect 14280 19508 14332 19514
rect 14280 19450 14332 19456
rect 14660 18426 14688 20402
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14200 17202 14320 17218
rect 14200 17196 14332 17202
rect 14200 17190 14280 17196
rect 14280 17138 14332 17144
rect 14096 15564 14148 15570
rect 14096 15506 14148 15512
rect 14004 13388 14056 13394
rect 14004 13330 14056 13336
rect 14016 12850 14044 13330
rect 14096 13320 14148 13326
rect 14096 13262 14148 13268
rect 14108 12918 14136 13262
rect 14096 12912 14148 12918
rect 14096 12854 14148 12860
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 14016 10674 14044 12786
rect 14278 12744 14334 12753
rect 14278 12679 14334 12688
rect 14292 12442 14320 12679
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14096 12164 14148 12170
rect 14096 12106 14148 12112
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14016 10130 14044 10610
rect 14108 10198 14136 12106
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14292 10606 14320 11086
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14292 10266 14320 10542
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14096 10192 14148 10198
rect 14096 10134 14148 10140
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 13924 8634 13952 9046
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 14016 8514 14044 10066
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 14108 8634 14136 9454
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 13924 8486 14044 8514
rect 13820 6384 13872 6390
rect 13820 6326 13872 6332
rect 13924 6118 13952 8486
rect 14292 6662 14320 10202
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14096 6316 14148 6322
rect 14096 6258 14148 6264
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13556 5030 13584 5102
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 13372 3126 13400 4422
rect 13556 3534 13584 4966
rect 13912 4820 13964 4826
rect 13912 4762 13964 4768
rect 13924 4146 13952 4762
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 14016 4078 14044 5170
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 13636 4004 13688 4010
rect 13636 3946 13688 3952
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13360 3120 13412 3126
rect 13360 3062 13412 3068
rect 13556 3058 13584 3470
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 13648 2774 13676 3946
rect 13832 3398 13860 4014
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 14108 2774 14136 6258
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 14200 4758 14228 6122
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 14188 4752 14240 4758
rect 14188 4694 14240 4700
rect 14292 4690 14320 4966
rect 14280 4684 14332 4690
rect 14280 4626 14332 4632
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14200 3738 14228 4558
rect 14292 4214 14320 4626
rect 14280 4208 14332 4214
rect 14280 4150 14332 4156
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14384 3618 14412 18022
rect 14568 17882 14596 18226
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 14464 13456 14516 13462
rect 14464 13398 14516 13404
rect 14476 12374 14504 13398
rect 14464 12368 14516 12374
rect 14568 12345 14596 17070
rect 14752 16726 14780 18022
rect 14740 16720 14792 16726
rect 14740 16662 14792 16668
rect 14844 14618 14872 27338
rect 14936 25362 14964 28018
rect 15028 28014 15056 28698
rect 15016 28008 15068 28014
rect 15016 27950 15068 27956
rect 15304 27402 15332 39238
rect 15488 39098 15516 39306
rect 15476 39092 15528 39098
rect 15476 39034 15528 39040
rect 15672 39030 15700 39442
rect 15844 39432 15896 39438
rect 15844 39374 15896 39380
rect 15660 39024 15712 39030
rect 15660 38966 15712 38972
rect 15856 37924 15884 39374
rect 15948 39098 15976 39442
rect 15936 39092 15988 39098
rect 15936 39034 15988 39040
rect 15936 38956 15988 38962
rect 15936 38898 15988 38904
rect 15948 38554 15976 38898
rect 16040 38894 16068 41386
rect 16224 41206 16252 42094
rect 16212 41200 16264 41206
rect 16212 41142 16264 41148
rect 16224 40610 16252 41142
rect 16316 40730 16344 42230
rect 16684 41818 16712 43250
rect 16776 42906 16804 43250
rect 16764 42900 16816 42906
rect 16764 42842 16816 42848
rect 16672 41812 16724 41818
rect 16672 41754 16724 41760
rect 16868 41414 16896 44474
rect 16776 41386 16896 41414
rect 16486 40896 16542 40905
rect 16486 40831 16542 40840
rect 16394 40760 16450 40769
rect 16304 40724 16356 40730
rect 16394 40695 16450 40704
rect 16304 40666 16356 40672
rect 16408 40662 16436 40695
rect 16132 40582 16252 40610
rect 16396 40656 16448 40662
rect 16396 40598 16448 40604
rect 16028 38888 16080 38894
rect 16028 38830 16080 38836
rect 15936 38548 15988 38554
rect 15936 38490 15988 38496
rect 15856 37896 15976 37924
rect 15660 37392 15712 37398
rect 15660 37334 15712 37340
rect 15568 37120 15620 37126
rect 15568 37062 15620 37068
rect 15580 36786 15608 37062
rect 15568 36780 15620 36786
rect 15568 36722 15620 36728
rect 15568 36100 15620 36106
rect 15568 36042 15620 36048
rect 15476 35692 15528 35698
rect 15476 35634 15528 35640
rect 15488 35562 15516 35634
rect 15476 35556 15528 35562
rect 15476 35498 15528 35504
rect 15384 35080 15436 35086
rect 15384 35022 15436 35028
rect 15396 33590 15424 35022
rect 15476 34196 15528 34202
rect 15476 34138 15528 34144
rect 15384 33584 15436 33590
rect 15384 33526 15436 33532
rect 15396 32570 15424 33526
rect 15384 32564 15436 32570
rect 15384 32506 15436 32512
rect 15384 32224 15436 32230
rect 15384 32166 15436 32172
rect 15292 27396 15344 27402
rect 15292 27338 15344 27344
rect 15292 27124 15344 27130
rect 15292 27066 15344 27072
rect 15108 26920 15160 26926
rect 15108 26862 15160 26868
rect 15120 26466 15148 26862
rect 15120 26450 15240 26466
rect 15120 26444 15252 26450
rect 15120 26438 15200 26444
rect 15200 26386 15252 26392
rect 15304 26314 15332 27066
rect 15292 26308 15344 26314
rect 15292 26250 15344 26256
rect 15292 25900 15344 25906
rect 15292 25842 15344 25848
rect 14924 25356 14976 25362
rect 14924 25298 14976 25304
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 14922 21584 14978 21593
rect 14922 21519 14924 21528
rect 14976 21519 14978 21528
rect 14924 21490 14976 21496
rect 15212 21486 15240 21830
rect 15200 21480 15252 21486
rect 15200 21422 15252 21428
rect 15304 20602 15332 25842
rect 15396 22094 15424 32166
rect 15488 29238 15516 34138
rect 15580 33930 15608 36042
rect 15672 35562 15700 37334
rect 15752 37256 15804 37262
rect 15752 37198 15804 37204
rect 15764 35834 15792 37198
rect 15844 36576 15896 36582
rect 15844 36518 15896 36524
rect 15752 35828 15804 35834
rect 15752 35770 15804 35776
rect 15856 35698 15884 36518
rect 15752 35692 15804 35698
rect 15752 35634 15804 35640
rect 15844 35692 15896 35698
rect 15844 35634 15896 35640
rect 15660 35556 15712 35562
rect 15660 35498 15712 35504
rect 15672 35170 15700 35498
rect 15764 35290 15792 35634
rect 15752 35284 15804 35290
rect 15752 35226 15804 35232
rect 15672 35142 15792 35170
rect 15660 34944 15712 34950
rect 15660 34886 15712 34892
rect 15568 33924 15620 33930
rect 15568 33866 15620 33872
rect 15580 33046 15608 33866
rect 15568 33040 15620 33046
rect 15568 32982 15620 32988
rect 15672 32910 15700 34886
rect 15660 32904 15712 32910
rect 15660 32846 15712 32852
rect 15660 32496 15712 32502
rect 15660 32438 15712 32444
rect 15568 32292 15620 32298
rect 15568 32234 15620 32240
rect 15580 31822 15608 32234
rect 15568 31816 15620 31822
rect 15568 31758 15620 31764
rect 15476 29232 15528 29238
rect 15476 29174 15528 29180
rect 15476 28960 15528 28966
rect 15476 28902 15528 28908
rect 15488 28626 15516 28902
rect 15476 28620 15528 28626
rect 15476 28562 15528 28568
rect 15476 28484 15528 28490
rect 15476 28426 15528 28432
rect 15488 28218 15516 28426
rect 15476 28212 15528 28218
rect 15476 28154 15528 28160
rect 15476 27396 15528 27402
rect 15476 27338 15528 27344
rect 15488 27130 15516 27338
rect 15476 27124 15528 27130
rect 15476 27066 15528 27072
rect 15580 24206 15608 31758
rect 15672 31142 15700 32438
rect 15660 31136 15712 31142
rect 15660 31078 15712 31084
rect 15672 30258 15700 31078
rect 15660 30252 15712 30258
rect 15660 30194 15712 30200
rect 15764 29850 15792 35142
rect 15844 33516 15896 33522
rect 15844 33458 15896 33464
rect 15752 29844 15804 29850
rect 15752 29786 15804 29792
rect 15856 29306 15884 33458
rect 15844 29300 15896 29306
rect 15844 29242 15896 29248
rect 15752 29232 15804 29238
rect 15752 29174 15804 29180
rect 15568 24200 15620 24206
rect 15568 24142 15620 24148
rect 15396 22066 15516 22094
rect 15384 21004 15436 21010
rect 15384 20946 15436 20952
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 14922 20496 14978 20505
rect 15396 20482 15424 20946
rect 15120 20466 15424 20482
rect 14922 20431 14924 20440
rect 14976 20431 14978 20440
rect 15108 20460 15424 20466
rect 14924 20402 14976 20408
rect 15160 20454 15424 20460
rect 15108 20402 15160 20408
rect 15290 20360 15346 20369
rect 15290 20295 15346 20304
rect 15200 19848 15252 19854
rect 15120 19796 15200 19802
rect 15120 19790 15252 19796
rect 15120 19774 15240 19790
rect 15016 18692 15068 18698
rect 15016 18634 15068 18640
rect 14924 18420 14976 18426
rect 14924 18362 14976 18368
rect 14936 18154 14964 18362
rect 15028 18290 15056 18634
rect 15016 18284 15068 18290
rect 15016 18226 15068 18232
rect 15120 18154 15148 19774
rect 15200 19712 15252 19718
rect 15200 19654 15252 19660
rect 15212 19446 15240 19654
rect 15200 19440 15252 19446
rect 15200 19382 15252 19388
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 15212 18358 15240 19110
rect 15200 18352 15252 18358
rect 15200 18294 15252 18300
rect 14924 18148 14976 18154
rect 14924 18090 14976 18096
rect 15108 18148 15160 18154
rect 15108 18090 15160 18096
rect 15016 17604 15068 17610
rect 15016 17546 15068 17552
rect 15028 17338 15056 17546
rect 15016 17332 15068 17338
rect 15016 17274 15068 17280
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 14924 16992 14976 16998
rect 14924 16934 14976 16940
rect 14936 16182 14964 16934
rect 15028 16794 15056 17138
rect 15016 16788 15068 16794
rect 15016 16730 15068 16736
rect 15120 16674 15148 18090
rect 15304 17814 15332 20295
rect 15292 17808 15344 17814
rect 15292 17750 15344 17756
rect 15396 17524 15424 20454
rect 15488 17678 15516 22066
rect 15660 22024 15712 22030
rect 15660 21966 15712 21972
rect 15568 21956 15620 21962
rect 15568 21898 15620 21904
rect 15580 21690 15608 21898
rect 15672 21690 15700 21966
rect 15568 21684 15620 21690
rect 15568 21626 15620 21632
rect 15660 21684 15712 21690
rect 15660 21626 15712 21632
rect 15764 21554 15792 29174
rect 15856 28558 15884 29242
rect 15948 28994 15976 37896
rect 16026 37360 16082 37369
rect 16026 37295 16028 37304
rect 16080 37295 16082 37304
rect 16028 37266 16080 37272
rect 16028 36712 16080 36718
rect 16028 36654 16080 36660
rect 16040 36174 16068 36654
rect 16028 36168 16080 36174
rect 16028 36110 16080 36116
rect 16040 30274 16068 36110
rect 16132 30938 16160 40582
rect 16500 40526 16528 40831
rect 16776 40526 16804 41386
rect 16856 41268 16908 41274
rect 16856 41210 16908 41216
rect 16488 40520 16540 40526
rect 16488 40462 16540 40468
rect 16764 40520 16816 40526
rect 16764 40462 16816 40468
rect 16868 40390 16896 41210
rect 17040 41200 17092 41206
rect 17040 41142 17092 41148
rect 17052 40730 17080 41142
rect 17040 40724 17092 40730
rect 17040 40666 17092 40672
rect 16948 40588 17000 40594
rect 16948 40530 17000 40536
rect 16580 40384 16632 40390
rect 16580 40326 16632 40332
rect 16856 40384 16908 40390
rect 16856 40326 16908 40332
rect 16304 39908 16356 39914
rect 16304 39850 16356 39856
rect 16212 38004 16264 38010
rect 16212 37946 16264 37952
rect 16224 36854 16252 37946
rect 16212 36848 16264 36854
rect 16212 36790 16264 36796
rect 16224 36378 16252 36790
rect 16212 36372 16264 36378
rect 16212 36314 16264 36320
rect 16212 35148 16264 35154
rect 16212 35090 16264 35096
rect 16224 33454 16252 35090
rect 16212 33448 16264 33454
rect 16212 33390 16264 33396
rect 16120 30932 16172 30938
rect 16120 30874 16172 30880
rect 16212 30592 16264 30598
rect 16212 30534 16264 30540
rect 16224 30394 16252 30534
rect 16212 30388 16264 30394
rect 16212 30330 16264 30336
rect 16040 30246 16252 30274
rect 15948 28966 16068 28994
rect 16040 28937 16068 28966
rect 16026 28928 16082 28937
rect 16026 28863 16082 28872
rect 16120 28756 16172 28762
rect 16120 28698 16172 28704
rect 15844 28552 15896 28558
rect 15844 28494 15896 28500
rect 16132 28082 16160 28698
rect 16120 28076 16172 28082
rect 16120 28018 16172 28024
rect 15844 27328 15896 27334
rect 15844 27270 15896 27276
rect 15856 26994 15884 27270
rect 15844 26988 15896 26994
rect 15844 26930 15896 26936
rect 16224 24138 16252 30246
rect 16316 30054 16344 39850
rect 16396 38888 16448 38894
rect 16396 38830 16448 38836
rect 16304 30048 16356 30054
rect 16304 29990 16356 29996
rect 16304 28008 16356 28014
rect 16304 27950 16356 27956
rect 16316 26042 16344 27950
rect 16304 26036 16356 26042
rect 16304 25978 16356 25984
rect 16212 24132 16264 24138
rect 16212 24074 16264 24080
rect 16224 23594 16252 24074
rect 16212 23588 16264 23594
rect 16212 23530 16264 23536
rect 16408 23118 16436 38830
rect 16488 38276 16540 38282
rect 16488 38218 16540 38224
rect 16500 38010 16528 38218
rect 16488 38004 16540 38010
rect 16488 37946 16540 37952
rect 16592 37398 16620 40326
rect 16960 40118 16988 40530
rect 16948 40112 17000 40118
rect 16948 40054 17000 40060
rect 16764 39636 16816 39642
rect 16764 39578 16816 39584
rect 16776 39284 16804 39578
rect 16684 39256 16804 39284
rect 16684 37618 16712 39256
rect 16960 38434 16988 40054
rect 16868 38418 16988 38434
rect 16856 38412 16988 38418
rect 16908 38406 16988 38412
rect 16856 38354 16908 38360
rect 16948 38344 17000 38350
rect 16948 38286 17000 38292
rect 17040 38344 17092 38350
rect 17040 38286 17092 38292
rect 16764 38276 16816 38282
rect 16764 38218 16816 38224
rect 16776 37806 16804 38218
rect 16856 38208 16908 38214
rect 16856 38150 16908 38156
rect 16764 37800 16816 37806
rect 16764 37742 16816 37748
rect 16684 37590 16804 37618
rect 16580 37392 16632 37398
rect 16580 37334 16632 37340
rect 16672 37188 16724 37194
rect 16672 37130 16724 37136
rect 16684 36922 16712 37130
rect 16672 36916 16724 36922
rect 16672 36858 16724 36864
rect 16672 35828 16724 35834
rect 16672 35770 16724 35776
rect 16684 35698 16712 35770
rect 16672 35692 16724 35698
rect 16672 35634 16724 35640
rect 16488 35216 16540 35222
rect 16488 35158 16540 35164
rect 16500 34678 16528 35158
rect 16488 34672 16540 34678
rect 16488 34614 16540 34620
rect 16672 34400 16724 34406
rect 16672 34342 16724 34348
rect 16684 34134 16712 34342
rect 16672 34128 16724 34134
rect 16672 34070 16724 34076
rect 16776 34066 16804 37590
rect 16868 37262 16896 38150
rect 16960 37466 16988 38286
rect 16948 37460 17000 37466
rect 16948 37402 17000 37408
rect 16856 37256 16908 37262
rect 16856 37198 16908 37204
rect 16960 36854 16988 37402
rect 16948 36848 17000 36854
rect 16948 36790 17000 36796
rect 16960 36378 16988 36790
rect 16948 36372 17000 36378
rect 16948 36314 17000 36320
rect 16948 35488 17000 35494
rect 16948 35430 17000 35436
rect 16856 34604 16908 34610
rect 16856 34546 16908 34552
rect 16868 34406 16896 34546
rect 16856 34400 16908 34406
rect 16856 34342 16908 34348
rect 16764 34060 16816 34066
rect 16764 34002 16816 34008
rect 16488 33992 16540 33998
rect 16488 33934 16540 33940
rect 16672 33992 16724 33998
rect 16672 33934 16724 33940
rect 16500 33658 16528 33934
rect 16684 33862 16712 33934
rect 16672 33856 16724 33862
rect 16672 33798 16724 33804
rect 16488 33652 16540 33658
rect 16488 33594 16540 33600
rect 16672 33448 16724 33454
rect 16672 33390 16724 33396
rect 16684 32366 16712 33390
rect 16776 33266 16804 34002
rect 16868 33454 16896 34342
rect 16960 33930 16988 35430
rect 16948 33924 17000 33930
rect 16948 33866 17000 33872
rect 16948 33584 17000 33590
rect 16948 33526 17000 33532
rect 16856 33448 16908 33454
rect 16856 33390 16908 33396
rect 16776 33238 16896 33266
rect 16764 32428 16816 32434
rect 16764 32370 16816 32376
rect 16672 32360 16724 32366
rect 16672 32302 16724 32308
rect 16672 32224 16724 32230
rect 16672 32166 16724 32172
rect 16488 31408 16540 31414
rect 16488 31350 16540 31356
rect 16500 30190 16528 31350
rect 16684 30784 16712 32166
rect 16776 31958 16804 32370
rect 16764 31952 16816 31958
rect 16764 31894 16816 31900
rect 16868 31754 16896 33238
rect 16592 30756 16712 30784
rect 16776 31726 16896 31754
rect 16488 30184 16540 30190
rect 16488 30126 16540 30132
rect 16120 23112 16172 23118
rect 16120 23054 16172 23060
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 15752 21548 15804 21554
rect 15752 21490 15804 21496
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15568 21412 15620 21418
rect 15568 21354 15620 21360
rect 15580 20466 15608 21354
rect 15660 20596 15712 20602
rect 15660 20538 15712 20544
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15580 20369 15608 20402
rect 15566 20360 15622 20369
rect 15566 20295 15622 20304
rect 15568 19984 15620 19990
rect 15568 19926 15620 19932
rect 15580 18902 15608 19926
rect 15568 18896 15620 18902
rect 15568 18838 15620 18844
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 15396 17496 15608 17524
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15028 16646 15148 16674
rect 15290 16688 15346 16697
rect 14924 16176 14976 16182
rect 14924 16118 14976 16124
rect 14924 15496 14976 15502
rect 15028 15484 15056 16646
rect 15290 16623 15346 16632
rect 15304 16590 15332 16623
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 15120 15706 15148 16526
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15108 15700 15160 15706
rect 15108 15642 15160 15648
rect 14976 15456 15056 15484
rect 14924 15438 14976 15444
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 15212 14482 15240 14758
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 15120 13938 15148 14214
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15120 13802 15148 13874
rect 15108 13796 15160 13802
rect 15108 13738 15160 13744
rect 15120 13326 15148 13738
rect 15212 13530 15240 14418
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 15304 13258 15332 15846
rect 15396 15706 15424 17138
rect 15488 16454 15516 17138
rect 15580 17134 15608 17496
rect 15568 17128 15620 17134
rect 15568 17070 15620 17076
rect 15580 16726 15608 17070
rect 15568 16720 15620 16726
rect 15568 16662 15620 16668
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 15672 15042 15700 20538
rect 15764 18902 15792 21490
rect 15856 21010 15884 21490
rect 15844 21004 15896 21010
rect 15844 20946 15896 20952
rect 16028 20256 16080 20262
rect 16028 20198 16080 20204
rect 16040 19378 16068 20198
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 15752 18896 15804 18902
rect 15752 18838 15804 18844
rect 15752 18760 15804 18766
rect 15752 18702 15804 18708
rect 15764 18086 15792 18702
rect 15948 18306 15976 19314
rect 15948 18290 16068 18306
rect 15948 18284 16080 18290
rect 15948 18278 16028 18284
rect 16028 18226 16080 18232
rect 15752 18080 15804 18086
rect 15752 18022 15804 18028
rect 16040 17610 16068 18226
rect 16028 17604 16080 17610
rect 16028 17546 16080 17552
rect 16040 17270 16068 17546
rect 15752 17264 15804 17270
rect 15752 17206 15804 17212
rect 16028 17264 16080 17270
rect 16028 17206 16080 17212
rect 15764 17066 15792 17206
rect 15936 17196 15988 17202
rect 15936 17138 15988 17144
rect 15752 17060 15804 17066
rect 15752 17002 15804 17008
rect 15764 16590 15792 17002
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15948 16250 15976 17138
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 16040 15502 16068 16934
rect 16028 15496 16080 15502
rect 16028 15438 16080 15444
rect 16132 15348 16160 23054
rect 16212 21956 16264 21962
rect 16212 21898 16264 21904
rect 16224 21146 16252 21898
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 16212 21140 16264 21146
rect 16212 21082 16264 21088
rect 16316 19854 16344 21830
rect 16488 21616 16540 21622
rect 16486 21584 16488 21593
rect 16540 21584 16542 21593
rect 16486 21519 16542 21528
rect 16500 20466 16528 21519
rect 16592 20874 16620 30756
rect 16672 30660 16724 30666
rect 16672 30602 16724 30608
rect 16684 30326 16712 30602
rect 16672 30320 16724 30326
rect 16672 30262 16724 30268
rect 16776 28506 16804 31726
rect 16856 31340 16908 31346
rect 16856 31282 16908 31288
rect 16868 30598 16896 31282
rect 16856 30592 16908 30598
rect 16856 30534 16908 30540
rect 16960 30410 16988 33526
rect 16684 28478 16804 28506
rect 16868 30382 16988 30410
rect 16684 27946 16712 28478
rect 16764 28416 16816 28422
rect 16764 28358 16816 28364
rect 16776 28150 16804 28358
rect 16764 28144 16816 28150
rect 16764 28086 16816 28092
rect 16672 27940 16724 27946
rect 16672 27882 16724 27888
rect 16764 27600 16816 27606
rect 16764 27542 16816 27548
rect 16776 27130 16804 27542
rect 16764 27124 16816 27130
rect 16764 27066 16816 27072
rect 16764 26784 16816 26790
rect 16764 26726 16816 26732
rect 16672 25968 16724 25974
rect 16672 25910 16724 25916
rect 16684 25226 16712 25910
rect 16672 25220 16724 25226
rect 16672 25162 16724 25168
rect 16684 24886 16712 25162
rect 16672 24880 16724 24886
rect 16672 24822 16724 24828
rect 16684 23050 16712 24822
rect 16776 24750 16804 26726
rect 16868 24818 16896 30382
rect 16948 30252 17000 30258
rect 16948 30194 17000 30200
rect 16960 30054 16988 30194
rect 16948 30048 17000 30054
rect 16948 29990 17000 29996
rect 16960 26042 16988 29990
rect 16948 26036 17000 26042
rect 16948 25978 17000 25984
rect 17052 25294 17080 38286
rect 17144 35834 17172 45902
rect 17224 45892 17276 45898
rect 17224 45834 17276 45840
rect 17236 43654 17264 45834
rect 17512 45490 17540 47738
rect 17880 47240 17908 49200
rect 17960 47252 18012 47258
rect 17880 47212 17960 47240
rect 17960 47194 18012 47200
rect 18144 47048 18196 47054
rect 18144 46990 18196 46996
rect 18236 47048 18288 47054
rect 18236 46990 18288 46996
rect 18052 46912 18104 46918
rect 18052 46854 18104 46860
rect 17868 46572 17920 46578
rect 17868 46514 17920 46520
rect 17776 46504 17828 46510
rect 17776 46446 17828 46452
rect 17500 45484 17552 45490
rect 17500 45426 17552 45432
rect 17316 45416 17368 45422
rect 17316 45358 17368 45364
rect 17328 44538 17356 45358
rect 17512 45014 17540 45426
rect 17500 45008 17552 45014
rect 17500 44950 17552 44956
rect 17316 44532 17368 44538
rect 17316 44474 17368 44480
rect 17500 43784 17552 43790
rect 17500 43726 17552 43732
rect 17224 43648 17276 43654
rect 17224 43590 17276 43596
rect 17236 40390 17264 43590
rect 17408 42628 17460 42634
rect 17408 42570 17460 42576
rect 17316 42084 17368 42090
rect 17316 42026 17368 42032
rect 17328 41002 17356 42026
rect 17316 40996 17368 41002
rect 17316 40938 17368 40944
rect 17316 40520 17368 40526
rect 17316 40462 17368 40468
rect 17224 40384 17276 40390
rect 17224 40326 17276 40332
rect 17224 40044 17276 40050
rect 17224 39986 17276 39992
rect 17236 39302 17264 39986
rect 17328 39982 17356 40462
rect 17316 39976 17368 39982
rect 17316 39918 17368 39924
rect 17224 39296 17276 39302
rect 17224 39238 17276 39244
rect 17236 38554 17264 39238
rect 17316 39024 17368 39030
rect 17316 38966 17368 38972
rect 17224 38548 17276 38554
rect 17224 38490 17276 38496
rect 17328 38418 17356 38966
rect 17316 38412 17368 38418
rect 17316 38354 17368 38360
rect 17420 38350 17448 42570
rect 17512 42362 17540 43726
rect 17500 42356 17552 42362
rect 17500 42298 17552 42304
rect 17684 41812 17736 41818
rect 17684 41754 17736 41760
rect 17696 41138 17724 41754
rect 17684 41132 17736 41138
rect 17684 41074 17736 41080
rect 17592 40996 17644 41002
rect 17592 40938 17644 40944
rect 17604 40458 17632 40938
rect 17592 40452 17644 40458
rect 17592 40394 17644 40400
rect 17592 38956 17644 38962
rect 17592 38898 17644 38904
rect 17604 38554 17632 38898
rect 17684 38752 17736 38758
rect 17684 38694 17736 38700
rect 17696 38554 17724 38694
rect 17592 38548 17644 38554
rect 17592 38490 17644 38496
rect 17684 38548 17736 38554
rect 17684 38490 17736 38496
rect 17408 38344 17460 38350
rect 17408 38286 17460 38292
rect 17682 37360 17738 37369
rect 17682 37295 17684 37304
rect 17736 37295 17738 37304
rect 17684 37266 17736 37272
rect 17788 37097 17816 46446
rect 17880 46102 17908 46514
rect 17868 46096 17920 46102
rect 17868 46038 17920 46044
rect 18064 44402 18092 46854
rect 18156 46170 18184 46990
rect 18248 46714 18276 46990
rect 18708 46918 18736 49200
rect 19536 47258 19564 49200
rect 20260 47932 20312 47938
rect 20260 47874 20312 47880
rect 19984 47592 20036 47598
rect 19984 47534 20036 47540
rect 19524 47252 19576 47258
rect 19524 47194 19576 47200
rect 19340 47048 19392 47054
rect 19340 46990 19392 46996
rect 18696 46912 18748 46918
rect 18696 46854 18748 46860
rect 19352 46714 19380 46990
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 18236 46708 18288 46714
rect 18236 46650 18288 46656
rect 19340 46708 19392 46714
rect 19340 46650 19392 46656
rect 18696 46572 18748 46578
rect 18696 46514 18748 46520
rect 18144 46164 18196 46170
rect 18144 46106 18196 46112
rect 18144 45620 18196 45626
rect 18144 45562 18196 45568
rect 18156 44878 18184 45562
rect 18708 45558 18736 46514
rect 19340 46504 19392 46510
rect 19340 46446 19392 46452
rect 18696 45552 18748 45558
rect 18696 45494 18748 45500
rect 18328 45484 18380 45490
rect 18328 45426 18380 45432
rect 18144 44872 18196 44878
rect 18144 44814 18196 44820
rect 18340 44538 18368 45426
rect 19352 45354 19380 46446
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19996 45490 20024 47534
rect 19984 45484 20036 45490
rect 19984 45426 20036 45432
rect 19340 45348 19392 45354
rect 19340 45290 19392 45296
rect 19996 44946 20024 45426
rect 18696 44940 18748 44946
rect 18696 44882 18748 44888
rect 19984 44940 20036 44946
rect 19984 44882 20036 44888
rect 18328 44532 18380 44538
rect 18328 44474 18380 44480
rect 18052 44396 18104 44402
rect 18052 44338 18104 44344
rect 18064 43858 18092 44338
rect 18144 44260 18196 44266
rect 18144 44202 18196 44208
rect 18052 43852 18104 43858
rect 18052 43794 18104 43800
rect 18156 43110 18184 44202
rect 18144 43104 18196 43110
rect 18144 43046 18196 43052
rect 18052 42220 18104 42226
rect 18052 42162 18104 42168
rect 17960 42016 18012 42022
rect 17960 41958 18012 41964
rect 17972 41206 18000 41958
rect 18064 41274 18092 42162
rect 18052 41268 18104 41274
rect 18052 41210 18104 41216
rect 17960 41200 18012 41206
rect 17960 41142 18012 41148
rect 17960 40520 18012 40526
rect 17960 40462 18012 40468
rect 17868 40180 17920 40186
rect 17868 40122 17920 40128
rect 17880 39370 17908 40122
rect 17972 39982 18000 40462
rect 17960 39976 18012 39982
rect 17960 39918 18012 39924
rect 17868 39364 17920 39370
rect 17868 39306 17920 39312
rect 17880 38282 17908 39306
rect 18156 39284 18184 43046
rect 18326 41304 18382 41313
rect 18326 41239 18328 41248
rect 18380 41239 18382 41248
rect 18328 41210 18380 41216
rect 18236 41200 18288 41206
rect 18234 41168 18236 41177
rect 18288 41168 18290 41177
rect 18234 41103 18290 41112
rect 18328 41132 18380 41138
rect 18328 41074 18380 41080
rect 18340 41041 18368 41074
rect 18326 41032 18382 41041
rect 18326 40967 18382 40976
rect 18328 40928 18380 40934
rect 18328 40870 18380 40876
rect 17972 39256 18184 39284
rect 18236 39296 18288 39302
rect 17868 38276 17920 38282
rect 17868 38218 17920 38224
rect 17880 37806 17908 38218
rect 17868 37800 17920 37806
rect 17868 37742 17920 37748
rect 17972 37262 18000 39256
rect 18236 39238 18288 39244
rect 18052 38548 18104 38554
rect 18052 38490 18104 38496
rect 18064 38350 18092 38490
rect 18248 38418 18276 39238
rect 18236 38412 18288 38418
rect 18236 38354 18288 38360
rect 18052 38344 18104 38350
rect 18052 38286 18104 38292
rect 18340 37874 18368 40870
rect 18512 40044 18564 40050
rect 18512 39986 18564 39992
rect 18524 39370 18552 39986
rect 18512 39364 18564 39370
rect 18512 39306 18564 39312
rect 18524 38758 18552 39306
rect 18512 38752 18564 38758
rect 18512 38694 18564 38700
rect 18420 38004 18472 38010
rect 18420 37946 18472 37952
rect 18432 37874 18460 37946
rect 18524 37942 18552 38694
rect 18512 37936 18564 37942
rect 18512 37878 18564 37884
rect 18328 37868 18380 37874
rect 18328 37810 18380 37816
rect 18420 37868 18472 37874
rect 18420 37810 18472 37816
rect 18604 37868 18656 37874
rect 18604 37810 18656 37816
rect 18236 37664 18288 37670
rect 18236 37606 18288 37612
rect 18248 37262 18276 37606
rect 17960 37256 18012 37262
rect 17960 37198 18012 37204
rect 18144 37256 18196 37262
rect 18144 37198 18196 37204
rect 18236 37256 18288 37262
rect 18236 37198 18288 37204
rect 17774 37088 17830 37097
rect 17774 37023 17830 37032
rect 17684 36780 17736 36786
rect 17684 36722 17736 36728
rect 17592 36712 17644 36718
rect 17592 36654 17644 36660
rect 17132 35828 17184 35834
rect 17132 35770 17184 35776
rect 17130 35728 17186 35737
rect 17130 35663 17186 35672
rect 17144 34610 17172 35663
rect 17132 34604 17184 34610
rect 17132 34546 17184 34552
rect 17144 33590 17172 34546
rect 17408 33992 17460 33998
rect 17408 33934 17460 33940
rect 17316 33856 17368 33862
rect 17316 33798 17368 33804
rect 17132 33584 17184 33590
rect 17132 33526 17184 33532
rect 17328 32434 17356 33798
rect 17420 32978 17448 33934
rect 17408 32972 17460 32978
rect 17408 32914 17460 32920
rect 17132 32428 17184 32434
rect 17132 32370 17184 32376
rect 17316 32428 17368 32434
rect 17316 32370 17368 32376
rect 17144 31346 17172 32370
rect 17316 32020 17368 32026
rect 17316 31962 17368 31968
rect 17132 31340 17184 31346
rect 17132 31282 17184 31288
rect 17132 31136 17184 31142
rect 17132 31078 17184 31084
rect 17224 31136 17276 31142
rect 17224 31078 17276 31084
rect 17144 30258 17172 31078
rect 17236 30394 17264 31078
rect 17328 30802 17356 31962
rect 17316 30796 17368 30802
rect 17316 30738 17368 30744
rect 17224 30388 17276 30394
rect 17224 30330 17276 30336
rect 17132 30252 17184 30258
rect 17132 30194 17184 30200
rect 17316 30252 17368 30258
rect 17316 30194 17368 30200
rect 17328 29646 17356 30194
rect 17316 29640 17368 29646
rect 17316 29582 17368 29588
rect 17420 29102 17448 32914
rect 17500 32224 17552 32230
rect 17500 32166 17552 32172
rect 17512 32026 17540 32166
rect 17500 32020 17552 32026
rect 17500 31962 17552 31968
rect 17604 31754 17632 36654
rect 17696 36174 17724 36722
rect 17788 36258 17816 37023
rect 17960 36712 18012 36718
rect 17960 36654 18012 36660
rect 17788 36230 17908 36258
rect 17684 36168 17736 36174
rect 17684 36110 17736 36116
rect 17696 35086 17724 36110
rect 17776 36100 17828 36106
rect 17776 36042 17828 36048
rect 17684 35080 17736 35086
rect 17684 35022 17736 35028
rect 17696 32774 17724 35022
rect 17788 34746 17816 36042
rect 17776 34740 17828 34746
rect 17776 34682 17828 34688
rect 17788 33454 17816 34682
rect 17880 34678 17908 36230
rect 17972 35290 18000 36654
rect 18156 36378 18184 37198
rect 18432 37194 18460 37810
rect 18512 37800 18564 37806
rect 18512 37742 18564 37748
rect 18328 37188 18380 37194
rect 18328 37130 18380 37136
rect 18420 37188 18472 37194
rect 18420 37130 18472 37136
rect 18340 36718 18368 37130
rect 18328 36712 18380 36718
rect 18328 36654 18380 36660
rect 18144 36372 18196 36378
rect 18144 36314 18196 36320
rect 18420 36236 18472 36242
rect 18420 36178 18472 36184
rect 17960 35284 18012 35290
rect 17960 35226 18012 35232
rect 18432 35086 18460 36178
rect 18420 35080 18472 35086
rect 18420 35022 18472 35028
rect 17868 34672 17920 34678
rect 17868 34614 17920 34620
rect 17960 34672 18012 34678
rect 17960 34614 18012 34620
rect 17972 34474 18000 34614
rect 18328 34604 18380 34610
rect 18328 34546 18380 34552
rect 17960 34468 18012 34474
rect 17960 34410 18012 34416
rect 17972 33998 18000 34410
rect 18236 34128 18288 34134
rect 18236 34070 18288 34076
rect 17960 33992 18012 33998
rect 17960 33934 18012 33940
rect 17868 33924 17920 33930
rect 17868 33866 17920 33872
rect 17880 33658 17908 33866
rect 17868 33652 17920 33658
rect 17868 33594 17920 33600
rect 17776 33448 17828 33454
rect 17776 33390 17828 33396
rect 17684 32768 17736 32774
rect 17684 32710 17736 32716
rect 17788 31754 17816 33390
rect 17880 32978 17908 33594
rect 17868 32972 17920 32978
rect 17868 32914 17920 32920
rect 17880 32502 17908 32914
rect 17868 32496 17920 32502
rect 17868 32438 17920 32444
rect 17868 32360 17920 32366
rect 17868 32302 17920 32308
rect 17512 31726 17632 31754
rect 17776 31748 17828 31754
rect 17408 29096 17460 29102
rect 17408 29038 17460 29044
rect 17512 28994 17540 31726
rect 17776 31690 17828 31696
rect 17776 30660 17828 30666
rect 17776 30602 17828 30608
rect 17788 30394 17816 30602
rect 17776 30388 17828 30394
rect 17776 30330 17828 30336
rect 17776 29164 17828 29170
rect 17696 29124 17776 29152
rect 17592 29096 17644 29102
rect 17592 29038 17644 29044
rect 17420 28966 17540 28994
rect 17420 27606 17448 28966
rect 17500 28076 17552 28082
rect 17500 28018 17552 28024
rect 17512 27674 17540 28018
rect 17500 27668 17552 27674
rect 17500 27610 17552 27616
rect 17408 27600 17460 27606
rect 17408 27542 17460 27548
rect 17222 27160 17278 27169
rect 17222 27095 17224 27104
rect 17276 27095 17278 27104
rect 17224 27066 17276 27072
rect 17316 25968 17368 25974
rect 17316 25910 17368 25916
rect 17040 25288 17092 25294
rect 17040 25230 17092 25236
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 16764 24744 16816 24750
rect 16764 24686 16816 24692
rect 16868 24614 16896 24754
rect 16856 24608 16908 24614
rect 16856 24550 16908 24556
rect 16672 23044 16724 23050
rect 16672 22986 16724 22992
rect 17052 22094 17080 25230
rect 17132 24812 17184 24818
rect 17132 24754 17184 24760
rect 17144 23866 17172 24754
rect 17328 24682 17356 25910
rect 17408 25900 17460 25906
rect 17408 25842 17460 25848
rect 17420 25498 17448 25842
rect 17408 25492 17460 25498
rect 17408 25434 17460 25440
rect 17604 25378 17632 29038
rect 17420 25350 17632 25378
rect 17316 24676 17368 24682
rect 17316 24618 17368 24624
rect 17328 24138 17356 24618
rect 17316 24132 17368 24138
rect 17316 24074 17368 24080
rect 17132 23860 17184 23866
rect 17132 23802 17184 23808
rect 17328 23798 17356 24074
rect 17316 23792 17368 23798
rect 17316 23734 17368 23740
rect 17224 23248 17276 23254
rect 17224 23190 17276 23196
rect 17236 23118 17264 23190
rect 17224 23112 17276 23118
rect 17224 23054 17276 23060
rect 16960 22066 17080 22094
rect 16856 21888 16908 21894
rect 16856 21830 16908 21836
rect 16764 21480 16816 21486
rect 16764 21422 16816 21428
rect 16776 20942 16804 21422
rect 16672 20936 16724 20942
rect 16672 20878 16724 20884
rect 16764 20936 16816 20942
rect 16764 20878 16816 20884
rect 16580 20868 16632 20874
rect 16580 20810 16632 20816
rect 16684 20482 16712 20878
rect 16868 20534 16896 21830
rect 16488 20460 16540 20466
rect 16488 20402 16540 20408
rect 16592 20454 16712 20482
rect 16856 20528 16908 20534
rect 16856 20470 16908 20476
rect 16764 20460 16816 20466
rect 16592 20262 16620 20454
rect 16764 20402 16816 20408
rect 16672 20324 16724 20330
rect 16672 20266 16724 20272
rect 16580 20256 16632 20262
rect 16580 20198 16632 20204
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 16396 19780 16448 19786
rect 16396 19722 16448 19728
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 16224 17542 16252 18702
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 16212 17536 16264 17542
rect 16212 17478 16264 17484
rect 16224 16697 16252 17478
rect 16210 16688 16266 16697
rect 16210 16623 16266 16632
rect 16212 16448 16264 16454
rect 16212 16390 16264 16396
rect 15580 15014 15700 15042
rect 16040 15320 16160 15348
rect 15476 14816 15528 14822
rect 15396 14764 15476 14770
rect 15396 14758 15528 14764
rect 15396 14742 15516 14758
rect 15396 14414 15424 14742
rect 15580 14550 15608 15014
rect 15660 14952 15712 14958
rect 15660 14894 15712 14900
rect 15568 14544 15620 14550
rect 15568 14486 15620 14492
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 15396 14074 15424 14350
rect 15672 14346 15700 14894
rect 15660 14340 15712 14346
rect 15660 14282 15712 14288
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 15672 14006 15700 14282
rect 15660 14000 15712 14006
rect 15660 13942 15712 13948
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15488 13734 15516 13874
rect 15568 13864 15620 13870
rect 15568 13806 15620 13812
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15488 13326 15516 13670
rect 15580 13326 15608 13806
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 15292 13252 15344 13258
rect 15292 13194 15344 13200
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15212 12434 15240 12786
rect 15212 12406 15424 12434
rect 14464 12310 14516 12316
rect 14554 12336 14610 12345
rect 14554 12271 14610 12280
rect 15014 12336 15070 12345
rect 15014 12271 15070 12280
rect 15028 10742 15056 12271
rect 15108 12232 15160 12238
rect 15108 12174 15160 12180
rect 15016 10736 15068 10742
rect 15016 10678 15068 10684
rect 15028 9926 15056 10678
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14844 8090 14872 8910
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14936 7886 14964 8230
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 14556 7812 14608 7818
rect 14556 7754 14608 7760
rect 14568 6458 14596 7754
rect 15120 6458 15148 12174
rect 15396 12170 15424 12406
rect 15488 12306 15516 13262
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15384 12164 15436 12170
rect 15384 12106 15436 12112
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 15212 10606 15240 11018
rect 15304 10674 15332 11086
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 15212 10266 15240 10542
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 15108 6452 15160 6458
rect 15108 6394 15160 6400
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14660 5846 14688 6054
rect 14648 5840 14700 5846
rect 14648 5782 14700 5788
rect 14648 5704 14700 5710
rect 14648 5646 14700 5652
rect 14660 5166 14688 5646
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14646 4312 14702 4321
rect 14646 4247 14702 4256
rect 14660 4146 14688 4247
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 12728 2746 12940 2774
rect 13004 2746 13124 2774
rect 13556 2746 13676 2774
rect 13924 2746 14136 2774
rect 14200 3590 14412 3618
rect 12728 800 12756 2746
rect 13004 2446 13032 2746
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 13096 800 13124 2246
rect 13556 800 13584 2746
rect 13924 800 13952 2746
rect 14200 2446 14228 3590
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 14292 800 14320 3130
rect 14476 3126 14504 3878
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 14476 2446 14504 3062
rect 14660 2854 14688 3334
rect 14648 2848 14700 2854
rect 14648 2790 14700 2796
rect 14660 2446 14688 2790
rect 14464 2440 14516 2446
rect 14464 2382 14516 2388
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 14752 1034 14780 6190
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14844 2650 14872 3470
rect 14936 2922 14964 4014
rect 14924 2916 14976 2922
rect 14924 2858 14976 2864
rect 14832 2644 14884 2650
rect 14832 2586 14884 2592
rect 14936 2514 14964 2858
rect 14924 2508 14976 2514
rect 14924 2450 14976 2456
rect 14660 1006 14780 1034
rect 14660 800 14688 1006
rect 15028 800 15056 6258
rect 15212 4282 15240 9930
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 15304 7750 15332 8230
rect 15396 7868 15424 12106
rect 15580 11218 15608 13262
rect 15672 12646 15700 13942
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15764 11626 15792 12378
rect 15752 11620 15804 11626
rect 15752 11562 15804 11568
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15488 8498 15516 8774
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15580 8022 15608 11018
rect 15672 10674 15700 11154
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15764 9654 15792 11562
rect 15856 11354 15884 13874
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15948 12714 15976 13262
rect 15936 12708 15988 12714
rect 15936 12650 15988 12656
rect 16040 12434 16068 15320
rect 16224 14482 16252 16390
rect 16212 14476 16264 14482
rect 16212 14418 16264 14424
rect 16120 13252 16172 13258
rect 16120 13194 16172 13200
rect 15948 12406 16068 12434
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 15752 9648 15804 9654
rect 15752 9590 15804 9596
rect 15660 9444 15712 9450
rect 15660 9386 15712 9392
rect 15672 8090 15700 9386
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15568 8016 15620 8022
rect 15568 7958 15620 7964
rect 15856 7954 15884 8366
rect 15948 8362 15976 12406
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 16040 11082 16068 12174
rect 16132 11694 16160 13194
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 16028 11076 16080 11082
rect 16028 11018 16080 11024
rect 16040 9994 16068 11018
rect 16132 10062 16160 11630
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 16028 9988 16080 9994
rect 16028 9930 16080 9936
rect 16028 9444 16080 9450
rect 16028 9386 16080 9392
rect 16040 9178 16068 9386
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 16132 8566 16160 9998
rect 16224 9178 16252 10610
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16224 8634 16252 9114
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16120 8560 16172 8566
rect 16120 8502 16172 8508
rect 15936 8356 15988 8362
rect 15936 8298 15988 8304
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 15476 7880 15528 7886
rect 15396 7840 15476 7868
rect 15476 7822 15528 7828
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15488 7546 15516 7822
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 16132 6866 16160 8502
rect 16224 7954 16252 8570
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 15476 6792 15528 6798
rect 16316 6746 16344 18566
rect 16408 18358 16436 19722
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 16592 18834 16620 19654
rect 16684 19242 16712 20266
rect 16776 19786 16804 20402
rect 16764 19780 16816 19786
rect 16764 19722 16816 19728
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16672 19236 16724 19242
rect 16672 19178 16724 19184
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 16580 18624 16632 18630
rect 16580 18566 16632 18572
rect 16396 18352 16448 18358
rect 16396 18294 16448 18300
rect 16396 16448 16448 16454
rect 16396 16390 16448 16396
rect 16408 12918 16436 16390
rect 16488 14544 16540 14550
rect 16486 14512 16488 14521
rect 16540 14512 16542 14521
rect 16486 14447 16542 14456
rect 16396 12912 16448 12918
rect 16396 12854 16448 12860
rect 16396 12776 16448 12782
rect 16396 12718 16448 12724
rect 16408 12646 16436 12718
rect 16396 12640 16448 12646
rect 16396 12582 16448 12588
rect 16408 12442 16436 12582
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16488 12300 16540 12306
rect 16488 12242 16540 12248
rect 16396 12164 16448 12170
rect 16396 12106 16448 12112
rect 16408 11694 16436 12106
rect 16396 11688 16448 11694
rect 16396 11630 16448 11636
rect 16408 10810 16436 11630
rect 16500 11558 16528 12242
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16408 9994 16436 10406
rect 16500 10266 16528 11494
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16396 9988 16448 9994
rect 16396 9930 16448 9936
rect 15476 6734 15528 6740
rect 15488 6390 15516 6734
rect 15948 6718 16344 6746
rect 15476 6384 15528 6390
rect 15476 6326 15528 6332
rect 15752 5840 15804 5846
rect 15752 5782 15804 5788
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15488 4690 15516 5510
rect 15476 4684 15528 4690
rect 15476 4626 15528 4632
rect 15292 4548 15344 4554
rect 15292 4490 15344 4496
rect 15304 4282 15332 4490
rect 15200 4276 15252 4282
rect 15200 4218 15252 4224
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 15198 4040 15254 4049
rect 15198 3975 15254 3984
rect 15212 3058 15240 3975
rect 15488 3942 15516 4626
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 15304 2774 15332 3878
rect 15672 3738 15700 4082
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15304 2746 15424 2774
rect 15396 800 15424 2746
rect 15764 2378 15792 5782
rect 15844 3392 15896 3398
rect 15844 3334 15896 3340
rect 15752 2372 15804 2378
rect 15752 2314 15804 2320
rect 15856 1034 15884 3334
rect 15948 2038 15976 6718
rect 16120 5772 16172 5778
rect 16120 5714 16172 5720
rect 15936 2032 15988 2038
rect 15936 1974 15988 1980
rect 15764 1006 15884 1034
rect 15764 800 15792 1006
rect 16132 800 16160 5714
rect 16212 5636 16264 5642
rect 16212 5578 16264 5584
rect 16224 4690 16252 5578
rect 16304 5092 16356 5098
rect 16304 5034 16356 5040
rect 16212 4684 16264 4690
rect 16212 4626 16264 4632
rect 16316 4622 16344 5034
rect 16304 4616 16356 4622
rect 16304 4558 16356 4564
rect 16316 4214 16344 4558
rect 16304 4208 16356 4214
rect 16304 4150 16356 4156
rect 16408 4010 16436 9930
rect 16488 5568 16540 5574
rect 16488 5510 16540 5516
rect 16500 4554 16528 5510
rect 16488 4548 16540 4554
rect 16488 4490 16540 4496
rect 16396 4004 16448 4010
rect 16396 3946 16448 3952
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 16500 800 16528 2246
rect 16592 2106 16620 18566
rect 16776 15366 16804 19450
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 16868 17882 16896 18702
rect 16856 17876 16908 17882
rect 16856 17818 16908 17824
rect 16868 16590 16896 17818
rect 16856 16584 16908 16590
rect 16856 16526 16908 16532
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 16672 15088 16724 15094
rect 16672 15030 16724 15036
rect 16684 14414 16712 15030
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16672 14408 16724 14414
rect 16724 14368 16804 14396
rect 16672 14350 16724 14356
rect 16672 13456 16724 13462
rect 16672 13398 16724 13404
rect 16684 12850 16712 13398
rect 16776 13326 16804 14368
rect 16868 14346 16896 14758
rect 16856 14340 16908 14346
rect 16856 14282 16908 14288
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16684 10810 16712 12786
rect 16764 12708 16816 12714
rect 16764 12650 16816 12656
rect 16776 12442 16804 12650
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16776 11762 16804 12378
rect 16868 12374 16896 14282
rect 16960 13530 16988 22066
rect 17316 22024 17368 22030
rect 17316 21966 17368 21972
rect 17328 21554 17356 21966
rect 17316 21548 17368 21554
rect 17316 21490 17368 21496
rect 17132 21480 17184 21486
rect 17132 21422 17184 21428
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 17052 18766 17080 20198
rect 17144 19514 17172 21422
rect 17224 20800 17276 20806
rect 17224 20742 17276 20748
rect 17132 19508 17184 19514
rect 17132 19450 17184 19456
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 17236 18630 17264 20742
rect 17328 20058 17356 21490
rect 17316 20052 17368 20058
rect 17316 19994 17368 20000
rect 17328 19378 17356 19994
rect 17316 19372 17368 19378
rect 17316 19314 17368 19320
rect 17224 18624 17276 18630
rect 17224 18566 17276 18572
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17236 17610 17264 18226
rect 17224 17604 17276 17610
rect 17224 17546 17276 17552
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 17052 16590 17080 16934
rect 17144 16658 17172 17478
rect 17236 17134 17264 17546
rect 17224 17128 17276 17134
rect 17224 17070 17276 17076
rect 17132 16652 17184 16658
rect 17132 16594 17184 16600
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 17040 16448 17092 16454
rect 17040 16390 17092 16396
rect 17052 16114 17080 16390
rect 17328 16182 17356 19314
rect 17316 16176 17368 16182
rect 17316 16118 17368 16124
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 17328 14006 17356 16118
rect 17420 15042 17448 25350
rect 17500 23724 17552 23730
rect 17500 23666 17552 23672
rect 17512 23322 17540 23666
rect 17500 23316 17552 23322
rect 17500 23258 17552 23264
rect 17500 22432 17552 22438
rect 17500 22374 17552 22380
rect 17512 21944 17540 22374
rect 17512 21916 17632 21944
rect 17604 18970 17632 21916
rect 17592 18964 17644 18970
rect 17592 18906 17644 18912
rect 17592 18284 17644 18290
rect 17592 18226 17644 18232
rect 17604 18193 17632 18226
rect 17590 18184 17646 18193
rect 17590 18119 17646 18128
rect 17604 17678 17632 18119
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17592 16584 17644 16590
rect 17590 16552 17592 16561
rect 17644 16552 17646 16561
rect 17590 16487 17646 16496
rect 17420 15014 17632 15042
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 17420 14278 17448 14894
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17316 14000 17368 14006
rect 17316 13942 17368 13948
rect 17224 13932 17276 13938
rect 17144 13892 17224 13920
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 17144 13326 17172 13892
rect 17224 13874 17276 13880
rect 17420 13394 17448 14214
rect 17512 13870 17540 14350
rect 17500 13864 17552 13870
rect 17500 13806 17552 13812
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 17040 12912 17092 12918
rect 17040 12854 17092 12860
rect 16856 12368 16908 12374
rect 16856 12310 16908 12316
rect 16856 11824 16908 11830
rect 16856 11766 16908 11772
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16868 11286 16896 11766
rect 16856 11280 16908 11286
rect 16856 11222 16908 11228
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16776 9926 16804 10610
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 16960 8974 16988 9522
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 16672 8900 16724 8906
rect 16672 8842 16724 8848
rect 16684 8022 16712 8842
rect 16672 8016 16724 8022
rect 16672 7958 16724 7964
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16684 6254 16712 7142
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16868 6254 16896 6598
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16948 6180 17000 6186
rect 16948 6122 17000 6128
rect 16960 5914 16988 6122
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 16776 4078 16804 5646
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16868 4622 16896 5102
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 16764 4072 16816 4078
rect 16764 4014 16816 4020
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16684 3466 16712 3878
rect 16764 3732 16816 3738
rect 16764 3674 16816 3680
rect 16672 3460 16724 3466
rect 16672 3402 16724 3408
rect 16776 3058 16804 3674
rect 16868 3534 16896 4558
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 16960 3738 16988 4422
rect 17052 4321 17080 12854
rect 17144 11898 17172 13262
rect 17604 12918 17632 15014
rect 17696 12918 17724 29124
rect 17880 29152 17908 32302
rect 17972 32065 18000 33934
rect 18248 33862 18276 34070
rect 18236 33856 18288 33862
rect 18236 33798 18288 33804
rect 18248 33522 18276 33798
rect 18340 33658 18368 34546
rect 18328 33652 18380 33658
rect 18328 33594 18380 33600
rect 18144 33516 18196 33522
rect 18144 33458 18196 33464
rect 18236 33516 18288 33522
rect 18236 33458 18288 33464
rect 18052 33448 18104 33454
rect 18052 33390 18104 33396
rect 17958 32056 18014 32065
rect 17958 31991 18014 32000
rect 18064 31822 18092 33390
rect 18052 31816 18104 31822
rect 18052 31758 18104 31764
rect 17960 31748 18012 31754
rect 17960 31690 18012 31696
rect 17828 29124 17908 29152
rect 17776 29106 17828 29112
rect 17972 28626 18000 31690
rect 18156 31686 18184 33458
rect 18328 33108 18380 33114
rect 18328 33050 18380 33056
rect 18236 32836 18288 32842
rect 18236 32778 18288 32784
rect 18248 32230 18276 32778
rect 18236 32224 18288 32230
rect 18236 32166 18288 32172
rect 18234 32056 18290 32065
rect 18234 31991 18290 32000
rect 18248 31958 18276 31991
rect 18236 31952 18288 31958
rect 18236 31894 18288 31900
rect 18144 31680 18196 31686
rect 18144 31622 18196 31628
rect 18156 31498 18184 31622
rect 18064 31470 18184 31498
rect 18236 31476 18288 31482
rect 18064 28694 18092 31470
rect 18236 31418 18288 31424
rect 18144 31340 18196 31346
rect 18144 31282 18196 31288
rect 18052 28688 18104 28694
rect 18052 28630 18104 28636
rect 17960 28620 18012 28626
rect 17960 28562 18012 28568
rect 17972 28098 18000 28562
rect 18052 28552 18104 28558
rect 18052 28494 18104 28500
rect 18064 28218 18092 28494
rect 18052 28212 18104 28218
rect 18052 28154 18104 28160
rect 17972 28070 18092 28098
rect 17868 28008 17920 28014
rect 17868 27950 17920 27956
rect 17776 26784 17828 26790
rect 17776 26726 17828 26732
rect 17788 24818 17816 26726
rect 17880 25702 17908 27950
rect 17960 26988 18012 26994
rect 17960 26930 18012 26936
rect 17972 26382 18000 26930
rect 17960 26376 18012 26382
rect 17960 26318 18012 26324
rect 17868 25696 17920 25702
rect 17868 25638 17920 25644
rect 17960 25356 18012 25362
rect 17960 25298 18012 25304
rect 17972 25158 18000 25298
rect 17960 25152 18012 25158
rect 17960 25094 18012 25100
rect 17776 24812 17828 24818
rect 17776 24754 17828 24760
rect 17960 24812 18012 24818
rect 17960 24754 18012 24760
rect 17788 22506 17816 24754
rect 17972 24614 18000 24754
rect 17960 24608 18012 24614
rect 17960 24550 18012 24556
rect 17776 22500 17828 22506
rect 17776 22442 17828 22448
rect 17960 22092 18012 22098
rect 17960 22034 18012 22040
rect 17972 21894 18000 22034
rect 17960 21888 18012 21894
rect 17880 21836 17960 21842
rect 17880 21830 18012 21836
rect 17880 21814 18000 21830
rect 17776 20936 17828 20942
rect 17776 20878 17828 20884
rect 17788 20602 17816 20878
rect 17776 20596 17828 20602
rect 17776 20538 17828 20544
rect 17880 20482 17908 21814
rect 17788 20454 17908 20482
rect 17960 20460 18012 20466
rect 17788 15314 17816 20454
rect 17960 20402 18012 20408
rect 17972 19446 18000 20402
rect 17960 19440 18012 19446
rect 17960 19382 18012 19388
rect 17868 19372 17920 19378
rect 17868 19314 17920 19320
rect 17880 18426 17908 19314
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 17868 17196 17920 17202
rect 17868 17138 17920 17144
rect 17880 16182 17908 17138
rect 17972 16454 18000 19382
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 17868 16176 17920 16182
rect 17868 16118 17920 16124
rect 17880 15502 17908 16118
rect 17868 15496 17920 15502
rect 17868 15438 17920 15444
rect 17972 15434 18000 16390
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 17788 15286 18000 15314
rect 17868 14816 17920 14822
rect 17868 14758 17920 14764
rect 17880 14414 17908 14758
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17880 13870 17908 14350
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17788 13308 17816 13806
rect 17880 13462 17908 13806
rect 17972 13802 18000 15286
rect 18064 14074 18092 28070
rect 18156 22778 18184 31282
rect 18248 31278 18276 31418
rect 18236 31272 18288 31278
rect 18236 31214 18288 31220
rect 18248 30258 18276 31214
rect 18340 31210 18368 33050
rect 18328 31204 18380 31210
rect 18328 31146 18380 31152
rect 18328 30592 18380 30598
rect 18328 30534 18380 30540
rect 18236 30252 18288 30258
rect 18236 30194 18288 30200
rect 18340 30190 18368 30534
rect 18328 30184 18380 30190
rect 18328 30126 18380 30132
rect 18328 30048 18380 30054
rect 18328 29990 18380 29996
rect 18236 28484 18288 28490
rect 18236 28426 18288 28432
rect 18248 22930 18276 28426
rect 18340 25378 18368 29990
rect 18432 26042 18460 35022
rect 18524 31414 18552 37742
rect 18616 37466 18644 37810
rect 18604 37460 18656 37466
rect 18604 37402 18656 37408
rect 18616 37262 18644 37402
rect 18604 37256 18656 37262
rect 18604 37198 18656 37204
rect 18708 36922 18736 44882
rect 19248 44872 19300 44878
rect 19248 44814 19300 44820
rect 18788 40384 18840 40390
rect 18788 40326 18840 40332
rect 18696 36916 18748 36922
rect 18696 36858 18748 36864
rect 18604 34400 18656 34406
rect 18604 34342 18656 34348
rect 18616 33522 18644 34342
rect 18696 33652 18748 33658
rect 18696 33594 18748 33600
rect 18604 33516 18656 33522
rect 18604 33458 18656 33464
rect 18604 32904 18656 32910
rect 18604 32846 18656 32852
rect 18512 31408 18564 31414
rect 18512 31350 18564 31356
rect 18512 30388 18564 30394
rect 18512 30330 18564 30336
rect 18524 30258 18552 30330
rect 18512 30252 18564 30258
rect 18512 30194 18564 30200
rect 18512 29572 18564 29578
rect 18512 29514 18564 29520
rect 18524 29034 18552 29514
rect 18512 29028 18564 29034
rect 18512 28970 18564 28976
rect 18616 28422 18644 32846
rect 18708 31822 18736 33594
rect 18800 31890 18828 40326
rect 19260 40186 19288 44814
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 20076 44396 20128 44402
rect 20076 44338 20128 44344
rect 19800 44328 19852 44334
rect 19800 44270 19852 44276
rect 19812 43790 19840 44270
rect 19984 43988 20036 43994
rect 19984 43930 20036 43936
rect 19800 43784 19852 43790
rect 19800 43726 19852 43732
rect 19340 43716 19392 43722
rect 19340 43658 19392 43664
rect 19352 42362 19380 43658
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19892 43308 19944 43314
rect 19892 43250 19944 43256
rect 19904 42634 19932 43250
rect 19996 42702 20024 43930
rect 19984 42696 20036 42702
rect 19984 42638 20036 42644
rect 19892 42628 19944 42634
rect 19892 42570 19944 42576
rect 19432 42560 19484 42566
rect 19432 42502 19484 42508
rect 19340 42356 19392 42362
rect 19340 42298 19392 42304
rect 19444 42208 19472 42502
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 20088 42362 20116 44338
rect 20272 43926 20300 47874
rect 20536 47456 20588 47462
rect 20536 47398 20588 47404
rect 20260 43920 20312 43926
rect 20260 43862 20312 43868
rect 20260 42696 20312 42702
rect 20260 42638 20312 42644
rect 20076 42356 20128 42362
rect 20076 42298 20128 42304
rect 19524 42220 19576 42226
rect 19444 42180 19524 42208
rect 19524 42162 19576 42168
rect 20272 42106 20300 42638
rect 20444 42560 20496 42566
rect 20444 42502 20496 42508
rect 20352 42220 20404 42226
rect 20352 42162 20404 42168
rect 19984 42084 20036 42090
rect 19984 42026 20036 42032
rect 20180 42078 20300 42106
rect 19340 41472 19392 41478
rect 19340 41414 19392 41420
rect 19352 40526 19380 41414
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19524 41064 19576 41070
rect 19524 41006 19576 41012
rect 19536 40662 19564 41006
rect 19524 40656 19576 40662
rect 19524 40598 19576 40604
rect 19340 40520 19392 40526
rect 19340 40462 19392 40468
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19248 40180 19300 40186
rect 19248 40122 19300 40128
rect 19340 39908 19392 39914
rect 19340 39850 19392 39856
rect 19352 38350 19380 39850
rect 19432 39432 19484 39438
rect 19432 39374 19484 39380
rect 19444 38486 19472 39374
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19432 38480 19484 38486
rect 19432 38422 19484 38428
rect 18880 38344 18932 38350
rect 18880 38286 18932 38292
rect 19340 38344 19392 38350
rect 19340 38286 19392 38292
rect 18892 37670 18920 38286
rect 19352 38010 19380 38286
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19340 38004 19392 38010
rect 19340 37946 19392 37952
rect 19432 37800 19484 37806
rect 19432 37742 19484 37748
rect 18880 37664 18932 37670
rect 18880 37606 18932 37612
rect 19156 37120 19208 37126
rect 19156 37062 19208 37068
rect 19340 37120 19392 37126
rect 19340 37062 19392 37068
rect 19168 36854 19196 37062
rect 19156 36848 19208 36854
rect 19156 36790 19208 36796
rect 19168 36242 19196 36790
rect 19248 36644 19300 36650
rect 19248 36586 19300 36592
rect 19156 36236 19208 36242
rect 19156 36178 19208 36184
rect 19260 36174 19288 36586
rect 19248 36168 19300 36174
rect 19248 36110 19300 36116
rect 19156 35692 19208 35698
rect 19076 35652 19156 35680
rect 18880 35012 18932 35018
rect 19076 35000 19104 35652
rect 19156 35634 19208 35640
rect 19260 35290 19288 36110
rect 19248 35284 19300 35290
rect 19248 35226 19300 35232
rect 19156 35148 19208 35154
rect 19208 35108 19288 35136
rect 19156 35090 19208 35096
rect 19156 35012 19208 35018
rect 19076 34972 19156 35000
rect 18880 34954 18932 34960
rect 19156 34954 19208 34960
rect 18788 31884 18840 31890
rect 18788 31826 18840 31832
rect 18696 31816 18748 31822
rect 18696 31758 18748 31764
rect 18696 31408 18748 31414
rect 18696 31350 18748 31356
rect 18604 28416 18656 28422
rect 18604 28358 18656 28364
rect 18604 28076 18656 28082
rect 18604 28018 18656 28024
rect 18420 26036 18472 26042
rect 18420 25978 18472 25984
rect 18432 25498 18460 25978
rect 18420 25492 18472 25498
rect 18420 25434 18472 25440
rect 18340 25350 18552 25378
rect 18328 24268 18380 24274
rect 18328 24210 18380 24216
rect 18340 23118 18368 24210
rect 18328 23112 18380 23118
rect 18328 23054 18380 23060
rect 18248 22902 18368 22930
rect 18144 22772 18196 22778
rect 18144 22714 18196 22720
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 18144 22432 18196 22438
rect 18144 22374 18196 22380
rect 18156 20466 18184 22374
rect 18248 22234 18276 22578
rect 18236 22228 18288 22234
rect 18236 22170 18288 22176
rect 18236 20868 18288 20874
rect 18236 20810 18288 20816
rect 18248 20466 18276 20810
rect 18340 20806 18368 22902
rect 18420 21548 18472 21554
rect 18420 21490 18472 21496
rect 18432 21146 18460 21490
rect 18420 21140 18472 21146
rect 18420 21082 18472 21088
rect 18328 20800 18380 20806
rect 18328 20742 18380 20748
rect 18144 20460 18196 20466
rect 18144 20402 18196 20408
rect 18236 20460 18288 20466
rect 18236 20402 18288 20408
rect 18248 20346 18276 20402
rect 18156 20318 18276 20346
rect 18328 20392 18380 20398
rect 18328 20334 18380 20340
rect 18156 16726 18184 20318
rect 18340 19990 18368 20334
rect 18420 20256 18472 20262
rect 18420 20198 18472 20204
rect 18328 19984 18380 19990
rect 18328 19926 18380 19932
rect 18432 19854 18460 20198
rect 18236 19848 18288 19854
rect 18420 19848 18472 19854
rect 18288 19808 18368 19836
rect 18236 19790 18288 19796
rect 18236 19440 18288 19446
rect 18236 19382 18288 19388
rect 18144 16720 18196 16726
rect 18144 16662 18196 16668
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 18156 15706 18184 16526
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 17868 13456 17920 13462
rect 17868 13398 17920 13404
rect 17868 13320 17920 13326
rect 17788 13280 17868 13308
rect 17868 13262 17920 13268
rect 17592 12912 17644 12918
rect 17592 12854 17644 12860
rect 17684 12912 17736 12918
rect 17684 12854 17736 12860
rect 17696 12442 17724 12854
rect 17684 12436 17736 12442
rect 17684 12378 17736 12384
rect 17880 12374 17908 13262
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 17972 11778 18000 12174
rect 18064 11898 18092 12786
rect 18052 11892 18104 11898
rect 18052 11834 18104 11840
rect 17972 11750 18092 11778
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 17236 10198 17264 10746
rect 17592 10668 17644 10674
rect 17592 10610 17644 10616
rect 17224 10192 17276 10198
rect 17224 10134 17276 10140
rect 17236 7410 17264 10134
rect 17500 9988 17552 9994
rect 17500 9930 17552 9936
rect 17512 9722 17540 9930
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 17604 6458 17632 10610
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 17972 8634 18000 10202
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17132 6316 17184 6322
rect 17132 6258 17184 6264
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 17038 4312 17094 4321
rect 17038 4247 17094 4256
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 16856 2848 16908 2854
rect 16856 2790 16908 2796
rect 16868 2446 16896 2790
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 16580 2100 16632 2106
rect 16580 2042 16632 2048
rect 16960 1034 16988 3538
rect 17052 2650 17080 4082
rect 17144 3670 17172 6258
rect 17316 6248 17368 6254
rect 17316 6190 17368 6196
rect 17328 5710 17356 6190
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 17236 3942 17264 5170
rect 17316 5024 17368 5030
rect 17316 4966 17368 4972
rect 17328 4554 17356 4966
rect 17316 4548 17368 4554
rect 17316 4490 17368 4496
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 17420 2774 17448 6258
rect 17788 5914 17816 8434
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17972 7342 18000 7890
rect 18064 7750 18092 11750
rect 18156 11370 18184 14894
rect 18248 11558 18276 19382
rect 18340 18766 18368 19808
rect 18420 19790 18472 19796
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18326 18592 18382 18601
rect 18326 18527 18382 18536
rect 18340 15026 18368 18527
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18328 14612 18380 14618
rect 18328 14554 18380 14560
rect 18340 14521 18368 14554
rect 18326 14512 18382 14521
rect 18326 14447 18382 14456
rect 18328 12844 18380 12850
rect 18328 12786 18380 12792
rect 18340 12170 18368 12786
rect 18328 12164 18380 12170
rect 18328 12106 18380 12112
rect 18340 11762 18368 12106
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 18156 11342 18276 11370
rect 18340 11354 18368 11698
rect 18248 11286 18276 11342
rect 18328 11348 18380 11354
rect 18328 11290 18380 11296
rect 18236 11280 18288 11286
rect 18236 11222 18288 11228
rect 18144 11212 18196 11218
rect 18144 11154 18196 11160
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 18052 7404 18104 7410
rect 18052 7346 18104 7352
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 17972 6798 18000 7278
rect 18064 7002 18092 7346
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 18156 6866 18184 11154
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 18156 6474 18184 6802
rect 18248 6798 18276 11222
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 18340 7954 18368 8978
rect 18328 7948 18380 7954
rect 18328 7890 18380 7896
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18156 6446 18276 6474
rect 18144 6384 18196 6390
rect 18144 6326 18196 6332
rect 17776 5908 17828 5914
rect 17776 5850 17828 5856
rect 17960 5228 18012 5234
rect 17960 5170 18012 5176
rect 17776 5092 17828 5098
rect 17776 5034 17828 5040
rect 17592 4820 17644 4826
rect 17592 4762 17644 4768
rect 17604 4010 17632 4762
rect 17788 4282 17816 5034
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 17776 4276 17828 4282
rect 17776 4218 17828 4224
rect 17592 4004 17644 4010
rect 17592 3946 17644 3952
rect 17776 4004 17828 4010
rect 17776 3946 17828 3952
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17696 3126 17724 3878
rect 17788 3602 17816 3946
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 17880 3058 17908 4558
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 17236 2746 17448 2774
rect 17040 2644 17092 2650
rect 17040 2586 17092 2592
rect 16868 1006 16988 1034
rect 16868 800 16896 1006
rect 17236 800 17264 2746
rect 17592 2304 17644 2310
rect 17592 2246 17644 2252
rect 17604 800 17632 2246
rect 17972 800 18000 5170
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 18064 4146 18092 4966
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 18156 2378 18184 6326
rect 18248 6322 18276 6446
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 18432 5386 18460 19654
rect 18524 17218 18552 25350
rect 18616 23322 18644 28018
rect 18708 26994 18736 31350
rect 18788 30932 18840 30938
rect 18788 30874 18840 30880
rect 18800 30394 18828 30874
rect 18788 30388 18840 30394
rect 18788 30330 18840 30336
rect 18696 26988 18748 26994
rect 18696 26930 18748 26936
rect 18696 26376 18748 26382
rect 18696 26318 18748 26324
rect 18708 23526 18736 26318
rect 18788 25696 18840 25702
rect 18788 25638 18840 25644
rect 18800 25226 18828 25638
rect 18788 25220 18840 25226
rect 18788 25162 18840 25168
rect 18892 23594 18920 34954
rect 19168 34678 19196 34954
rect 18972 34672 19024 34678
rect 18972 34614 19024 34620
rect 19156 34672 19208 34678
rect 19156 34614 19208 34620
rect 19260 34626 19288 35108
rect 19352 34746 19380 37062
rect 19340 34740 19392 34746
rect 19340 34682 19392 34688
rect 18984 34474 19012 34614
rect 18972 34468 19024 34474
rect 18972 34410 19024 34416
rect 18984 33590 19012 34410
rect 19062 34096 19118 34105
rect 19062 34031 19118 34040
rect 19076 33930 19104 34031
rect 19064 33924 19116 33930
rect 19064 33866 19116 33872
rect 18972 33584 19024 33590
rect 18972 33526 19024 33532
rect 19168 30870 19196 34614
rect 19260 34598 19380 34626
rect 19352 34542 19380 34598
rect 19340 34536 19392 34542
rect 19340 34478 19392 34484
rect 19248 34400 19300 34406
rect 19248 34342 19300 34348
rect 19444 34354 19472 37742
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19892 36780 19944 36786
rect 19892 36722 19944 36728
rect 19616 36576 19668 36582
rect 19616 36518 19668 36524
rect 19628 36378 19656 36518
rect 19616 36372 19668 36378
rect 19616 36314 19668 36320
rect 19904 36310 19932 36722
rect 19892 36304 19944 36310
rect 19892 36246 19944 36252
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19708 35624 19760 35630
rect 19708 35566 19760 35572
rect 19720 35154 19748 35566
rect 19708 35148 19760 35154
rect 19708 35090 19760 35096
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19708 34672 19760 34678
rect 19708 34614 19760 34620
rect 19720 34474 19748 34614
rect 19708 34468 19760 34474
rect 19708 34410 19760 34416
rect 19260 33998 19288 34342
rect 19444 34326 19564 34354
rect 19432 34196 19484 34202
rect 19432 34138 19484 34144
rect 19444 33998 19472 34138
rect 19248 33992 19300 33998
rect 19248 33934 19300 33940
rect 19432 33992 19484 33998
rect 19432 33934 19484 33940
rect 19536 33912 19564 34326
rect 19996 33946 20024 42026
rect 20076 39296 20128 39302
rect 20076 39238 20128 39244
rect 20088 38962 20116 39238
rect 20076 38956 20128 38962
rect 20076 38898 20128 38904
rect 20076 38276 20128 38282
rect 20076 38218 20128 38224
rect 20088 38010 20116 38218
rect 20076 38004 20128 38010
rect 20076 37946 20128 37952
rect 20180 37126 20208 42078
rect 20260 42016 20312 42022
rect 20260 41958 20312 41964
rect 20272 40390 20300 41958
rect 20260 40384 20312 40390
rect 20260 40326 20312 40332
rect 20272 40118 20300 40326
rect 20260 40112 20312 40118
rect 20260 40054 20312 40060
rect 20260 39840 20312 39846
rect 20260 39782 20312 39788
rect 20272 38554 20300 39782
rect 20260 38548 20312 38554
rect 20260 38490 20312 38496
rect 20168 37120 20220 37126
rect 20168 37062 20220 37068
rect 20364 36632 20392 42162
rect 20456 42022 20484 42502
rect 20444 42016 20496 42022
rect 20444 41958 20496 41964
rect 20444 40996 20496 41002
rect 20444 40938 20496 40944
rect 20272 36604 20392 36632
rect 20168 36576 20220 36582
rect 20168 36518 20220 36524
rect 20076 35692 20128 35698
rect 20076 35634 20128 35640
rect 20088 34513 20116 35634
rect 20074 34504 20130 34513
rect 20074 34439 20130 34448
rect 20074 34096 20130 34105
rect 20074 34031 20076 34040
rect 20128 34031 20130 34040
rect 20076 34002 20128 34008
rect 19624 33924 19676 33930
rect 19536 33884 19624 33912
rect 19536 33844 19564 33884
rect 19996 33918 20116 33946
rect 19624 33866 19676 33872
rect 19516 33816 19564 33844
rect 19984 33856 20036 33862
rect 19516 33640 19544 33816
rect 19984 33798 20036 33804
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19516 33612 19564 33640
rect 19340 33108 19392 33114
rect 19340 33050 19392 33056
rect 19248 32904 19300 32910
rect 19248 32846 19300 32852
rect 19260 32502 19288 32846
rect 19248 32496 19300 32502
rect 19248 32438 19300 32444
rect 19352 31822 19380 33050
rect 19536 32910 19564 33612
rect 19432 32904 19484 32910
rect 19432 32846 19484 32852
rect 19524 32904 19576 32910
rect 19708 32904 19760 32910
rect 19524 32846 19576 32852
rect 19706 32872 19708 32881
rect 19760 32872 19762 32881
rect 19444 32026 19472 32846
rect 19536 32756 19564 32846
rect 19706 32807 19762 32816
rect 19516 32728 19564 32756
rect 19516 32552 19544 32728
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19516 32524 19564 32552
rect 19536 32298 19564 32524
rect 19524 32292 19576 32298
rect 19524 32234 19576 32240
rect 19432 32020 19484 32026
rect 19432 31962 19484 31968
rect 19340 31816 19392 31822
rect 19340 31758 19392 31764
rect 19156 30864 19208 30870
rect 19156 30806 19208 30812
rect 19352 30682 19380 31758
rect 19996 31754 20024 33798
rect 20088 33114 20116 33918
rect 20076 33108 20128 33114
rect 20076 33050 20128 33056
rect 19432 31748 19484 31754
rect 19996 31726 20116 31754
rect 19432 31690 19484 31696
rect 19444 31414 19472 31690
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19432 31408 19484 31414
rect 19432 31350 19484 31356
rect 19524 30864 19576 30870
rect 19524 30806 19576 30812
rect 19984 30864 20036 30870
rect 19984 30806 20036 30812
rect 19352 30654 19472 30682
rect 19536 30666 19564 30806
rect 19340 30592 19392 30598
rect 19340 30534 19392 30540
rect 19352 30326 19380 30534
rect 19340 30320 19392 30326
rect 19340 30262 19392 30268
rect 19444 30054 19472 30654
rect 19524 30660 19576 30666
rect 19524 30602 19576 30608
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19432 30048 19484 30054
rect 19432 29990 19484 29996
rect 19524 30048 19576 30054
rect 19524 29990 19576 29996
rect 19430 29880 19486 29889
rect 19430 29815 19486 29824
rect 19248 29572 19300 29578
rect 19248 29514 19300 29520
rect 19340 29572 19392 29578
rect 19340 29514 19392 29520
rect 19064 28416 19116 28422
rect 19064 28358 19116 28364
rect 19076 28218 19104 28358
rect 19064 28212 19116 28218
rect 19064 28154 19116 28160
rect 19076 27674 19104 28154
rect 19260 27946 19288 29514
rect 19248 27940 19300 27946
rect 19248 27882 19300 27888
rect 19352 27878 19380 29514
rect 19444 28422 19472 29815
rect 19536 29782 19564 29990
rect 19524 29776 19576 29782
rect 19524 29718 19576 29724
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19892 28960 19944 28966
rect 19892 28902 19944 28908
rect 19798 28656 19854 28665
rect 19798 28591 19800 28600
rect 19852 28591 19854 28600
rect 19800 28562 19852 28568
rect 19904 28558 19932 28902
rect 19524 28552 19576 28558
rect 19708 28552 19760 28558
rect 19524 28494 19576 28500
rect 19706 28520 19708 28529
rect 19892 28552 19944 28558
rect 19760 28520 19762 28529
rect 19432 28416 19484 28422
rect 19536 28404 19564 28494
rect 19892 28494 19944 28500
rect 19706 28455 19762 28464
rect 19432 28358 19484 28364
rect 19516 28376 19564 28404
rect 19516 28200 19544 28376
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19516 28172 19564 28200
rect 19432 28144 19484 28150
rect 19432 28086 19484 28092
rect 19340 27872 19392 27878
rect 19340 27814 19392 27820
rect 19338 27704 19394 27713
rect 19064 27668 19116 27674
rect 19338 27639 19394 27648
rect 19064 27610 19116 27616
rect 19352 27606 19380 27639
rect 19340 27600 19392 27606
rect 19340 27542 19392 27548
rect 19338 27432 19394 27441
rect 18972 27396 19024 27402
rect 19338 27367 19394 27376
rect 18972 27338 19024 27344
rect 18984 26450 19012 27338
rect 19248 27328 19300 27334
rect 19248 27270 19300 27276
rect 19260 26994 19288 27270
rect 19248 26988 19300 26994
rect 19248 26930 19300 26936
rect 18972 26444 19024 26450
rect 18972 26386 19024 26392
rect 18984 25974 19012 26386
rect 19352 26042 19380 27367
rect 19444 27062 19472 28086
rect 19536 27985 19564 28172
rect 19996 28150 20024 30806
rect 19984 28144 20036 28150
rect 19890 28112 19946 28121
rect 19984 28086 20036 28092
rect 19890 28047 19946 28056
rect 19522 27976 19578 27985
rect 19904 27946 19932 28047
rect 19522 27911 19578 27920
rect 19892 27940 19944 27946
rect 19892 27882 19944 27888
rect 19524 27872 19576 27878
rect 19524 27814 19576 27820
rect 19536 27470 19564 27814
rect 19892 27668 19944 27674
rect 19892 27610 19944 27616
rect 19708 27600 19760 27606
rect 19708 27542 19760 27548
rect 19720 27470 19748 27542
rect 19524 27464 19576 27470
rect 19524 27406 19576 27412
rect 19708 27464 19760 27470
rect 19904 27441 19932 27610
rect 19708 27406 19760 27412
rect 19890 27432 19946 27441
rect 19890 27367 19946 27376
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19432 27056 19484 27062
rect 19432 26998 19484 27004
rect 19340 26036 19392 26042
rect 19340 25978 19392 25984
rect 18972 25968 19024 25974
rect 18972 25910 19024 25916
rect 19340 25492 19392 25498
rect 19340 25434 19392 25440
rect 19064 24948 19116 24954
rect 19064 24890 19116 24896
rect 18972 24812 19024 24818
rect 18972 24754 19024 24760
rect 18984 24614 19012 24754
rect 18972 24608 19024 24614
rect 18972 24550 19024 24556
rect 18880 23588 18932 23594
rect 18880 23530 18932 23536
rect 18696 23520 18748 23526
rect 18696 23462 18748 23468
rect 18604 23316 18656 23322
rect 18604 23258 18656 23264
rect 18604 23112 18656 23118
rect 18604 23054 18656 23060
rect 18616 21690 18644 23054
rect 18708 21894 18736 23462
rect 18892 23254 18920 23530
rect 18880 23248 18932 23254
rect 18880 23190 18932 23196
rect 18984 23100 19012 24550
rect 18892 23072 19012 23100
rect 18788 22568 18840 22574
rect 18788 22510 18840 22516
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 18604 21684 18656 21690
rect 18604 21626 18656 21632
rect 18708 21554 18736 21830
rect 18800 21690 18828 22510
rect 18788 21684 18840 21690
rect 18788 21626 18840 21632
rect 18696 21548 18748 21554
rect 18696 21490 18748 21496
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18708 19938 18736 20742
rect 18800 20534 18828 21626
rect 18788 20528 18840 20534
rect 18788 20470 18840 20476
rect 18708 19910 18828 19938
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18708 18766 18736 19790
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18616 18290 18644 18702
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 18602 18184 18658 18193
rect 18602 18119 18604 18128
rect 18656 18119 18658 18128
rect 18604 18090 18656 18096
rect 18708 17338 18736 18702
rect 18696 17332 18748 17338
rect 18696 17274 18748 17280
rect 18524 17190 18736 17218
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18616 15706 18644 17070
rect 18604 15700 18656 15706
rect 18604 15642 18656 15648
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18616 12850 18644 14962
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18512 11552 18564 11558
rect 18512 11494 18564 11500
rect 18524 9674 18552 11494
rect 18616 11218 18644 12786
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18708 10266 18736 17190
rect 18800 13258 18828 19910
rect 18892 18737 18920 23072
rect 19076 22094 19104 24890
rect 19352 24750 19380 25434
rect 19444 24818 19472 26998
rect 19996 26994 20024 28086
rect 19984 26988 20036 26994
rect 19984 26930 20036 26936
rect 19984 26852 20036 26858
rect 19984 26794 20036 26800
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19996 25974 20024 26794
rect 19984 25968 20036 25974
rect 19984 25910 20036 25916
rect 19706 25392 19762 25401
rect 19706 25327 19708 25336
rect 19760 25327 19762 25336
rect 19708 25298 19760 25304
rect 19708 25220 19760 25226
rect 19760 25180 20024 25208
rect 19708 25162 19760 25168
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19996 24886 20024 25180
rect 19984 24880 20036 24886
rect 19984 24822 20036 24828
rect 19432 24812 19484 24818
rect 19432 24754 19484 24760
rect 19340 24744 19392 24750
rect 19340 24686 19392 24692
rect 19524 24608 19576 24614
rect 19576 24568 19748 24596
rect 19524 24550 19576 24556
rect 19522 24304 19578 24313
rect 19340 24268 19392 24274
rect 19522 24239 19578 24248
rect 19340 24210 19392 24216
rect 19352 24177 19380 24210
rect 19536 24206 19564 24239
rect 19720 24206 19748 24568
rect 19524 24200 19576 24206
rect 19338 24168 19394 24177
rect 19524 24142 19576 24148
rect 19708 24200 19760 24206
rect 19708 24142 19760 24148
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 19338 24103 19394 24112
rect 19294 24064 19346 24070
rect 19346 24012 19380 24018
rect 19294 24006 19380 24012
rect 19306 23990 19380 24006
rect 19352 23769 19380 23990
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19996 23798 20024 24142
rect 19524 23792 19576 23798
rect 19338 23760 19394 23769
rect 19338 23695 19394 23704
rect 19522 23760 19524 23769
rect 19984 23792 20036 23798
rect 19576 23760 19578 23769
rect 19984 23734 20036 23740
rect 19522 23695 19578 23704
rect 19154 23624 19210 23633
rect 19154 23559 19210 23568
rect 19168 23526 19196 23559
rect 19156 23520 19208 23526
rect 19156 23462 19208 23468
rect 20088 23066 20116 31726
rect 20180 27962 20208 36518
rect 20272 29578 20300 36604
rect 20352 35080 20404 35086
rect 20352 35022 20404 35028
rect 20364 34678 20392 35022
rect 20352 34672 20404 34678
rect 20456 34649 20484 40938
rect 20548 39914 20576 47398
rect 20640 47240 20668 49286
rect 21178 49200 21234 50000
rect 22006 49200 22062 50000
rect 22834 49314 22890 50000
rect 22834 49286 23152 49314
rect 22834 49200 22890 49286
rect 20720 47252 20772 47258
rect 20640 47212 20720 47240
rect 20720 47194 20772 47200
rect 21088 47184 21140 47190
rect 21088 47126 21140 47132
rect 20720 47048 20772 47054
rect 20720 46990 20772 46996
rect 20732 46714 20760 46990
rect 20720 46708 20772 46714
rect 20720 46650 20772 46656
rect 21100 45490 21128 47126
rect 21192 46696 21220 49200
rect 22020 47274 22048 49200
rect 22468 48000 22520 48006
rect 22468 47942 22520 47948
rect 22020 47258 22140 47274
rect 22020 47252 22152 47258
rect 22020 47246 22100 47252
rect 22100 47194 22152 47200
rect 22100 47048 22152 47054
rect 22100 46990 22152 46996
rect 22112 46714 22140 46990
rect 22100 46708 22152 46714
rect 21192 46668 21312 46696
rect 21180 46572 21232 46578
rect 21180 46514 21232 46520
rect 21192 45558 21220 46514
rect 21284 46442 21312 46668
rect 22100 46650 22152 46656
rect 21364 46640 21416 46646
rect 21364 46582 21416 46588
rect 21272 46436 21324 46442
rect 21272 46378 21324 46384
rect 21180 45552 21232 45558
rect 21180 45494 21232 45500
rect 21088 45484 21140 45490
rect 21008 45444 21088 45472
rect 20628 45416 20680 45422
rect 20628 45358 20680 45364
rect 20640 43994 20668 45358
rect 21008 44402 21036 45444
rect 21088 45426 21140 45432
rect 21088 45348 21140 45354
rect 21088 45290 21140 45296
rect 20996 44396 21048 44402
rect 20996 44338 21048 44344
rect 21100 44198 21128 45290
rect 21376 45082 21404 46582
rect 22376 45960 22428 45966
rect 22376 45902 22428 45908
rect 22388 45558 22416 45902
rect 22376 45552 22428 45558
rect 22376 45494 22428 45500
rect 22480 45490 22508 47942
rect 23124 47258 23152 49286
rect 23662 49200 23718 50000
rect 24490 49200 24546 50000
rect 25318 49200 25374 50000
rect 26146 49200 26202 50000
rect 27066 49200 27122 50000
rect 27894 49200 27950 50000
rect 28722 49314 28778 50000
rect 29550 49314 29606 50000
rect 28722 49286 28948 49314
rect 28722 49200 28778 49286
rect 23676 47258 23704 49200
rect 23112 47252 23164 47258
rect 23112 47194 23164 47200
rect 23664 47252 23716 47258
rect 23664 47194 23716 47200
rect 22928 47048 22980 47054
rect 22928 46990 22980 46996
rect 24400 47048 24452 47054
rect 24400 46990 24452 46996
rect 22940 46170 22968 46990
rect 23388 46980 23440 46986
rect 23388 46922 23440 46928
rect 23940 46980 23992 46986
rect 23940 46922 23992 46928
rect 22928 46164 22980 46170
rect 22928 46106 22980 46112
rect 23296 46028 23348 46034
rect 23296 45970 23348 45976
rect 23308 45626 23336 45970
rect 23296 45620 23348 45626
rect 23296 45562 23348 45568
rect 22468 45484 22520 45490
rect 22468 45426 22520 45432
rect 21364 45076 21416 45082
rect 21364 45018 21416 45024
rect 22480 44946 22508 45426
rect 22928 45416 22980 45422
rect 22928 45358 22980 45364
rect 22940 45286 22968 45358
rect 22928 45280 22980 45286
rect 22928 45222 22980 45228
rect 22468 44940 22520 44946
rect 22468 44882 22520 44888
rect 21732 44804 21784 44810
rect 21732 44746 21784 44752
rect 21088 44192 21140 44198
rect 21088 44134 21140 44140
rect 20628 43988 20680 43994
rect 20628 43930 20680 43936
rect 20720 43716 20772 43722
rect 20720 43658 20772 43664
rect 20628 43104 20680 43110
rect 20628 43046 20680 43052
rect 20640 42226 20668 43046
rect 20732 42838 20760 43658
rect 21100 43382 21128 44134
rect 21088 43376 21140 43382
rect 21088 43318 21140 43324
rect 20720 42832 20772 42838
rect 20720 42774 20772 42780
rect 20904 42832 20956 42838
rect 20904 42774 20956 42780
rect 20720 42628 20772 42634
rect 20720 42570 20772 42576
rect 20628 42220 20680 42226
rect 20628 42162 20680 42168
rect 20536 39908 20588 39914
rect 20536 39850 20588 39856
rect 20536 39296 20588 39302
rect 20536 39238 20588 39244
rect 20352 34614 20404 34620
rect 20442 34640 20498 34649
rect 20442 34575 20498 34584
rect 20352 34536 20404 34542
rect 20350 34504 20352 34513
rect 20404 34504 20406 34513
rect 20350 34439 20406 34448
rect 20364 33844 20392 34439
rect 20444 34400 20496 34406
rect 20444 34342 20496 34348
rect 20456 33998 20484 34342
rect 20548 34202 20576 39238
rect 20732 38350 20760 42570
rect 20916 42294 20944 42774
rect 20904 42288 20956 42294
rect 20904 42230 20956 42236
rect 20812 42220 20864 42226
rect 20812 42162 20864 42168
rect 20824 41070 20852 42162
rect 20916 41614 20944 42230
rect 20904 41608 20956 41614
rect 20904 41550 20956 41556
rect 20812 41064 20864 41070
rect 20812 41006 20864 41012
rect 20812 40520 20864 40526
rect 20812 40462 20864 40468
rect 20824 38554 20852 40462
rect 21100 39522 21128 43318
rect 21180 42696 21232 42702
rect 21180 42638 21232 42644
rect 21192 42226 21220 42638
rect 21180 42220 21232 42226
rect 21180 42162 21232 42168
rect 21456 42152 21508 42158
rect 21456 42094 21508 42100
rect 21180 41608 21232 41614
rect 21180 41550 21232 41556
rect 21192 40594 21220 41550
rect 21364 41064 21416 41070
rect 21364 41006 21416 41012
rect 21180 40588 21232 40594
rect 21180 40530 21232 40536
rect 21376 40526 21404 41006
rect 21468 40730 21496 42094
rect 21640 41200 21692 41206
rect 21640 41142 21692 41148
rect 21548 40928 21600 40934
rect 21548 40870 21600 40876
rect 21456 40724 21508 40730
rect 21456 40666 21508 40672
rect 21364 40520 21416 40526
rect 21364 40462 21416 40468
rect 21560 40118 21588 40870
rect 21652 40730 21680 41142
rect 21640 40724 21692 40730
rect 21640 40666 21692 40672
rect 21548 40112 21600 40118
rect 21548 40054 21600 40060
rect 20916 39494 21128 39522
rect 20812 38548 20864 38554
rect 20812 38490 20864 38496
rect 20720 38344 20772 38350
rect 20720 38286 20772 38292
rect 20628 37868 20680 37874
rect 20628 37810 20680 37816
rect 20812 37868 20864 37874
rect 20812 37810 20864 37816
rect 20640 36666 20668 37810
rect 20720 37120 20772 37126
rect 20720 37062 20772 37068
rect 20732 36786 20760 37062
rect 20720 36780 20772 36786
rect 20720 36722 20772 36728
rect 20640 36638 20760 36666
rect 20628 36100 20680 36106
rect 20628 36042 20680 36048
rect 20640 35630 20668 36042
rect 20628 35624 20680 35630
rect 20628 35566 20680 35572
rect 20628 35080 20680 35086
rect 20628 35022 20680 35028
rect 20536 34196 20588 34202
rect 20536 34138 20588 34144
rect 20534 34096 20590 34105
rect 20534 34031 20590 34040
rect 20548 33998 20576 34031
rect 20444 33992 20496 33998
rect 20444 33934 20496 33940
rect 20536 33992 20588 33998
rect 20536 33934 20588 33940
rect 20364 33816 20576 33844
rect 20444 33652 20496 33658
rect 20444 33594 20496 33600
rect 20456 33454 20484 33594
rect 20352 33448 20404 33454
rect 20352 33390 20404 33396
rect 20444 33448 20496 33454
rect 20444 33390 20496 33396
rect 20364 32774 20392 33390
rect 20548 33046 20576 33816
rect 20536 33040 20588 33046
rect 20536 32982 20588 32988
rect 20442 32872 20498 32881
rect 20442 32807 20498 32816
rect 20352 32768 20404 32774
rect 20352 32710 20404 32716
rect 20456 32570 20484 32807
rect 20444 32564 20496 32570
rect 20444 32506 20496 32512
rect 20352 32428 20404 32434
rect 20352 32370 20404 32376
rect 20364 31142 20392 32370
rect 20536 32360 20588 32366
rect 20536 32302 20588 32308
rect 20444 32292 20496 32298
rect 20444 32234 20496 32240
rect 20456 31822 20484 32234
rect 20548 31890 20576 32302
rect 20536 31884 20588 31890
rect 20536 31826 20588 31832
rect 20444 31816 20496 31822
rect 20444 31758 20496 31764
rect 20352 31136 20404 31142
rect 20352 31078 20404 31084
rect 20352 30252 20404 30258
rect 20352 30194 20404 30200
rect 20260 29572 20312 29578
rect 20260 29514 20312 29520
rect 20364 28642 20392 30194
rect 20536 29028 20588 29034
rect 20536 28970 20588 28976
rect 20444 28756 20496 28762
rect 20444 28698 20496 28704
rect 20272 28614 20392 28642
rect 20272 28082 20300 28614
rect 20456 28529 20484 28698
rect 20548 28558 20576 28970
rect 20536 28552 20588 28558
rect 20442 28520 20498 28529
rect 20536 28494 20588 28500
rect 20442 28455 20498 28464
rect 20534 28384 20590 28393
rect 20534 28319 20590 28328
rect 20260 28076 20312 28082
rect 20260 28018 20312 28024
rect 20180 27934 20392 27962
rect 20168 27872 20220 27878
rect 20168 27814 20220 27820
rect 19352 23038 20116 23066
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 19156 22228 19208 22234
rect 19156 22170 19208 22176
rect 18984 22066 19104 22094
rect 18984 19446 19012 22066
rect 19064 21956 19116 21962
rect 19064 21898 19116 21904
rect 19076 21690 19104 21898
rect 19064 21684 19116 21690
rect 19064 21626 19116 21632
rect 18972 19440 19024 19446
rect 18972 19382 19024 19388
rect 19076 18873 19104 21626
rect 19062 18864 19118 18873
rect 19062 18799 19118 18808
rect 18878 18728 18934 18737
rect 18878 18663 18934 18672
rect 19064 18624 19116 18630
rect 19064 18566 19116 18572
rect 18970 18456 19026 18465
rect 18970 18391 19026 18400
rect 18788 13252 18840 13258
rect 18788 13194 18840 13200
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 18892 12345 18920 12786
rect 18878 12336 18934 12345
rect 18878 12271 18934 12280
rect 18984 12102 19012 18391
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 18972 11756 19024 11762
rect 18972 11698 19024 11704
rect 18880 10736 18932 10742
rect 18880 10678 18932 10684
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18524 9646 18644 9674
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18524 8634 18552 8910
rect 18616 8838 18644 9646
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 18708 9178 18736 9522
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18616 8498 18644 8774
rect 18788 8560 18840 8566
rect 18788 8502 18840 8508
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18708 8362 18736 8434
rect 18696 8356 18748 8362
rect 18696 8298 18748 8304
rect 18512 8288 18564 8294
rect 18512 8230 18564 8236
rect 18524 7886 18552 8230
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18340 5358 18460 5386
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 18248 4214 18276 4422
rect 18236 4208 18288 4214
rect 18236 4150 18288 4156
rect 18248 4078 18276 4150
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 18340 3924 18368 5358
rect 18420 5228 18472 5234
rect 18420 5170 18472 5176
rect 18248 3896 18368 3924
rect 18248 2446 18276 3896
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 18340 3126 18368 3334
rect 18328 3120 18380 3126
rect 18328 3062 18380 3068
rect 18432 2774 18460 5170
rect 18524 4146 18552 7686
rect 18602 6896 18658 6905
rect 18602 6831 18658 6840
rect 18616 6458 18644 6831
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18708 6322 18736 6394
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18616 5642 18644 6190
rect 18708 6118 18736 6258
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 18604 5636 18656 5642
rect 18604 5578 18656 5584
rect 18800 5370 18828 8502
rect 18892 7954 18920 10678
rect 18880 7948 18932 7954
rect 18880 7890 18932 7896
rect 18880 6180 18932 6186
rect 18880 6122 18932 6128
rect 18892 5710 18920 6122
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18984 5574 19012 11698
rect 18972 5568 19024 5574
rect 18972 5510 19024 5516
rect 18788 5364 18840 5370
rect 18788 5306 18840 5312
rect 18972 5024 19024 5030
rect 18972 4966 19024 4972
rect 18984 4826 19012 4966
rect 18972 4820 19024 4826
rect 18972 4762 19024 4768
rect 19076 4434 19104 18566
rect 19168 14958 19196 22170
rect 19260 21622 19288 22578
rect 19248 21616 19300 21622
rect 19248 21558 19300 21564
rect 19260 20806 19288 21558
rect 19248 20800 19300 20806
rect 19248 20742 19300 20748
rect 19260 18902 19288 20742
rect 19248 18896 19300 18902
rect 19248 18838 19300 18844
rect 19352 18834 19380 23038
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19984 22772 20036 22778
rect 19984 22714 20036 22720
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19444 20806 19472 20878
rect 19432 20800 19484 20806
rect 19432 20742 19484 20748
rect 19444 19394 19472 20742
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19444 19366 19564 19394
rect 19432 19304 19484 19310
rect 19432 19246 19484 19252
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19352 18358 19380 18770
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 19444 17678 19472 19246
rect 19536 18737 19564 19366
rect 19996 19009 20024 22714
rect 20076 21956 20128 21962
rect 20076 21898 20128 21904
rect 20088 20602 20116 21898
rect 20076 20596 20128 20602
rect 20076 20538 20128 20544
rect 20074 20496 20130 20505
rect 20074 20431 20076 20440
rect 20128 20431 20130 20440
rect 20076 20402 20128 20408
rect 20180 20346 20208 27814
rect 20260 27464 20312 27470
rect 20260 27406 20312 27412
rect 20272 26790 20300 27406
rect 20260 26784 20312 26790
rect 20260 26726 20312 26732
rect 20260 25696 20312 25702
rect 20260 25638 20312 25644
rect 20272 25294 20300 25638
rect 20260 25288 20312 25294
rect 20260 25230 20312 25236
rect 20272 24206 20300 25230
rect 20260 24200 20312 24206
rect 20260 24142 20312 24148
rect 20258 23216 20314 23225
rect 20258 23151 20314 23160
rect 20272 23118 20300 23151
rect 20260 23112 20312 23118
rect 20260 23054 20312 23060
rect 20260 22976 20312 22982
rect 20260 22918 20312 22924
rect 20272 20466 20300 22918
rect 20260 20460 20312 20466
rect 20260 20402 20312 20408
rect 20076 20324 20128 20330
rect 20180 20318 20300 20346
rect 20076 20266 20128 20272
rect 19982 19000 20038 19009
rect 19982 18935 20038 18944
rect 19522 18728 19578 18737
rect 19522 18663 19578 18672
rect 19984 18692 20036 18698
rect 19984 18634 20036 18640
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19996 18442 20024 18634
rect 20088 18601 20116 20266
rect 20168 19780 20220 19786
rect 20168 19722 20220 19728
rect 20074 18592 20130 18601
rect 20074 18527 20130 18536
rect 19996 18414 20116 18442
rect 20180 18426 20208 19722
rect 19892 18284 19944 18290
rect 19892 18226 19944 18232
rect 19616 18216 19668 18222
rect 19616 18158 19668 18164
rect 19628 17882 19656 18158
rect 19708 18148 19760 18154
rect 19708 18090 19760 18096
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19720 17785 19748 18090
rect 19904 17921 19932 18226
rect 19982 18048 20038 18057
rect 19982 17983 20038 17992
rect 19890 17912 19946 17921
rect 19890 17847 19946 17856
rect 19706 17776 19762 17785
rect 19706 17711 19762 17720
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 19248 17060 19300 17066
rect 19248 17002 19300 17008
rect 19260 15994 19288 17002
rect 19352 16182 19380 17546
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19522 17232 19578 17241
rect 19522 17167 19524 17176
rect 19576 17167 19578 17176
rect 19524 17138 19576 17144
rect 19432 17128 19484 17134
rect 19432 17070 19484 17076
rect 19340 16176 19392 16182
rect 19340 16118 19392 16124
rect 19260 15966 19380 15994
rect 19352 14958 19380 15966
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19444 14822 19472 17070
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19706 15464 19762 15473
rect 19706 15399 19708 15408
rect 19760 15399 19762 15408
rect 19708 15370 19760 15376
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19340 14408 19392 14414
rect 19260 14356 19340 14362
rect 19260 14350 19392 14356
rect 19260 14334 19380 14350
rect 19432 14340 19484 14346
rect 19260 13818 19288 14334
rect 19432 14282 19484 14288
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19352 14006 19380 14214
rect 19340 14000 19392 14006
rect 19340 13942 19392 13948
rect 19260 13790 19380 13818
rect 19352 13462 19380 13790
rect 19340 13456 19392 13462
rect 19340 13398 19392 13404
rect 19444 13326 19472 14282
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19432 13320 19484 13326
rect 19352 13280 19432 13308
rect 19156 13252 19208 13258
rect 19156 13194 19208 13200
rect 19168 12850 19196 13194
rect 19352 12918 19380 13280
rect 19432 13262 19484 13268
rect 19432 13184 19484 13190
rect 19432 13126 19484 13132
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 19444 12850 19472 13126
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19996 12918 20024 17983
rect 20088 17678 20116 18414
rect 20168 18420 20220 18426
rect 20168 18362 20220 18368
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 20088 17338 20116 17614
rect 20076 17332 20128 17338
rect 20076 17274 20128 17280
rect 20166 17232 20222 17241
rect 20166 17167 20168 17176
rect 20220 17167 20222 17176
rect 20168 17138 20220 17144
rect 20074 17096 20130 17105
rect 20074 17031 20130 17040
rect 20168 17060 20220 17066
rect 20088 16998 20116 17031
rect 20168 17002 20220 17008
rect 20076 16992 20128 16998
rect 20076 16934 20128 16940
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 20088 16182 20116 16390
rect 20180 16250 20208 17002
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 20076 16176 20128 16182
rect 20076 16118 20128 16124
rect 20076 15972 20128 15978
rect 20076 15914 20128 15920
rect 20088 14618 20116 15914
rect 20166 15192 20222 15201
rect 20166 15127 20222 15136
rect 20180 15094 20208 15127
rect 20168 15088 20220 15094
rect 20168 15030 20220 15036
rect 20168 14816 20220 14822
rect 20168 14758 20220 14764
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 19984 12912 20036 12918
rect 19984 12854 20036 12860
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19444 12714 19472 12786
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 19798 12472 19854 12481
rect 19798 12407 19800 12416
rect 19852 12407 19854 12416
rect 19800 12378 19852 12384
rect 19248 12232 19300 12238
rect 20088 12186 20116 14350
rect 20180 13870 20208 14758
rect 20168 13864 20220 13870
rect 20168 13806 20220 13812
rect 19248 12174 19300 12180
rect 19260 11150 19288 12174
rect 19996 12158 20116 12186
rect 20166 12200 20222 12209
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19996 11898 20024 12158
rect 20166 12135 20222 12144
rect 20076 12096 20128 12102
rect 20076 12038 20128 12044
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 20088 11694 20116 12038
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 19432 11620 19484 11626
rect 19432 11562 19484 11568
rect 19708 11620 19760 11626
rect 19984 11620 20036 11626
rect 19760 11580 19840 11608
rect 19708 11562 19760 11568
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 19260 10010 19288 11086
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 19352 10606 19380 10950
rect 19444 10742 19472 11562
rect 19812 11150 19840 11580
rect 19984 11562 20036 11568
rect 19800 11144 19852 11150
rect 19800 11086 19852 11092
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19432 10736 19484 10742
rect 19432 10678 19484 10684
rect 19340 10600 19392 10606
rect 19340 10542 19392 10548
rect 19996 10470 20024 11562
rect 20076 11076 20128 11082
rect 20076 11018 20128 11024
rect 20088 10810 20116 11018
rect 20076 10804 20128 10810
rect 20076 10746 20128 10752
rect 20180 10690 20208 12135
rect 20272 11354 20300 20318
rect 20364 19938 20392 27934
rect 20444 27872 20496 27878
rect 20444 27814 20496 27820
rect 20456 24313 20484 27814
rect 20442 24304 20498 24313
rect 20442 24239 20498 24248
rect 20456 23594 20484 24239
rect 20444 23588 20496 23594
rect 20444 23530 20496 23536
rect 20548 21706 20576 28319
rect 20640 27878 20668 35022
rect 20732 34066 20760 36638
rect 20720 34060 20772 34066
rect 20720 34002 20772 34008
rect 20732 30274 20760 34002
rect 20824 31346 20852 37810
rect 20916 34746 20944 39494
rect 21088 39432 21140 39438
rect 21088 39374 21140 39380
rect 20996 39364 21048 39370
rect 20996 39306 21048 39312
rect 21008 38282 21036 39306
rect 21100 39098 21128 39374
rect 21456 39296 21508 39302
rect 21456 39238 21508 39244
rect 21088 39092 21140 39098
rect 21088 39034 21140 39040
rect 21180 38548 21232 38554
rect 21180 38490 21232 38496
rect 20996 38276 21048 38282
rect 20996 38218 21048 38224
rect 21008 37942 21036 38218
rect 21088 38208 21140 38214
rect 21088 38150 21140 38156
rect 21100 38010 21128 38150
rect 21088 38004 21140 38010
rect 21088 37946 21140 37952
rect 20996 37936 21048 37942
rect 20996 37878 21048 37884
rect 20996 37256 21048 37262
rect 20994 37224 20996 37233
rect 21048 37224 21050 37233
rect 20994 37159 21050 37168
rect 21088 37188 21140 37194
rect 21088 37130 21140 37136
rect 21100 36718 21128 37130
rect 20996 36712 21048 36718
rect 20996 36654 21048 36660
rect 21088 36712 21140 36718
rect 21088 36654 21140 36660
rect 21008 35494 21036 36654
rect 20996 35488 21048 35494
rect 20996 35430 21048 35436
rect 20996 35080 21048 35086
rect 20996 35022 21048 35028
rect 20904 34740 20956 34746
rect 20904 34682 20956 34688
rect 20904 34468 20956 34474
rect 20904 34410 20956 34416
rect 20916 33454 20944 34410
rect 21008 33522 21036 35022
rect 21088 33856 21140 33862
rect 21088 33798 21140 33804
rect 20996 33516 21048 33522
rect 20996 33458 21048 33464
rect 20904 33448 20956 33454
rect 20904 33390 20956 33396
rect 20904 31748 20956 31754
rect 20904 31690 20956 31696
rect 20916 31482 20944 31690
rect 20904 31476 20956 31482
rect 20904 31418 20956 31424
rect 20812 31340 20864 31346
rect 20812 31282 20864 31288
rect 20824 30394 20852 31282
rect 20812 30388 20864 30394
rect 20812 30330 20864 30336
rect 20732 30246 20944 30274
rect 20720 29232 20772 29238
rect 20720 29174 20772 29180
rect 20628 27872 20680 27878
rect 20628 27814 20680 27820
rect 20732 27690 20760 29174
rect 20812 29164 20864 29170
rect 20812 29106 20864 29112
rect 20824 28762 20852 29106
rect 20812 28756 20864 28762
rect 20812 28698 20864 28704
rect 20916 28608 20944 30246
rect 20640 27662 20760 27690
rect 20824 28580 20944 28608
rect 20640 27062 20668 27662
rect 20718 27568 20774 27577
rect 20718 27503 20774 27512
rect 20628 27056 20680 27062
rect 20628 26998 20680 27004
rect 20640 26450 20668 26998
rect 20628 26444 20680 26450
rect 20628 26386 20680 26392
rect 20628 25152 20680 25158
rect 20628 25094 20680 25100
rect 20640 24256 20668 25094
rect 20732 24954 20760 27503
rect 20824 26926 20852 28580
rect 20904 28484 20956 28490
rect 20904 28426 20956 28432
rect 20916 28218 20944 28426
rect 21008 28422 21036 33458
rect 20996 28416 21048 28422
rect 20996 28358 21048 28364
rect 20904 28212 20956 28218
rect 20904 28154 20956 28160
rect 20996 28076 21048 28082
rect 20996 28018 21048 28024
rect 20902 27976 20958 27985
rect 20902 27911 20958 27920
rect 20916 27878 20944 27911
rect 20904 27872 20956 27878
rect 20904 27814 20956 27820
rect 20916 27470 20944 27814
rect 21008 27674 21036 28018
rect 20996 27668 21048 27674
rect 20996 27610 21048 27616
rect 20904 27464 20956 27470
rect 20904 27406 20956 27412
rect 20812 26920 20864 26926
rect 20812 26862 20864 26868
rect 20904 26784 20956 26790
rect 20904 26726 20956 26732
rect 20916 26382 20944 26726
rect 20904 26376 20956 26382
rect 20904 26318 20956 26324
rect 20720 24948 20772 24954
rect 20720 24890 20772 24896
rect 20720 24268 20772 24274
rect 20640 24228 20720 24256
rect 20720 24210 20772 24216
rect 20626 24168 20682 24177
rect 20626 24103 20628 24112
rect 20680 24103 20682 24112
rect 20628 24074 20680 24080
rect 20732 23186 20760 24210
rect 20996 23656 21048 23662
rect 20996 23598 21048 23604
rect 20720 23180 20772 23186
rect 20720 23122 20772 23128
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 20720 22500 20772 22506
rect 20720 22442 20772 22448
rect 20732 22012 20760 22442
rect 20824 22166 20852 23054
rect 20904 23044 20956 23050
rect 20904 22986 20956 22992
rect 20916 22234 20944 22986
rect 20904 22228 20956 22234
rect 20904 22170 20956 22176
rect 20812 22160 20864 22166
rect 20812 22102 20864 22108
rect 20732 21984 20852 22012
rect 20548 21678 20760 21706
rect 20444 20460 20496 20466
rect 20444 20402 20496 20408
rect 20456 20097 20484 20402
rect 20442 20088 20498 20097
rect 20442 20023 20498 20032
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 20364 19910 20576 19938
rect 20444 19848 20496 19854
rect 20444 19790 20496 19796
rect 20456 19514 20484 19790
rect 20444 19508 20496 19514
rect 20444 19450 20496 19456
rect 20456 19378 20484 19450
rect 20444 19372 20496 19378
rect 20444 19314 20496 19320
rect 20352 18692 20404 18698
rect 20352 18634 20404 18640
rect 20364 18290 20392 18634
rect 20352 18284 20404 18290
rect 20352 18226 20404 18232
rect 20350 18048 20406 18057
rect 20350 17983 20406 17992
rect 20364 17626 20392 17983
rect 20456 17814 20484 19314
rect 20444 17808 20496 17814
rect 20444 17750 20496 17756
rect 20364 17598 20484 17626
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 20364 13954 20392 17478
rect 20456 15570 20484 17598
rect 20548 17270 20576 19910
rect 20536 17264 20588 17270
rect 20536 17206 20588 17212
rect 20536 16992 20588 16998
rect 20536 16934 20588 16940
rect 20548 16590 20576 16934
rect 20640 16590 20668 19994
rect 20732 18193 20760 21678
rect 20824 20058 20852 21984
rect 20904 21480 20956 21486
rect 20904 21422 20956 21428
rect 20916 20534 20944 21422
rect 20904 20528 20956 20534
rect 20904 20470 20956 20476
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 21008 19122 21036 23598
rect 21100 20262 21128 33798
rect 21192 31754 21220 38490
rect 21468 38350 21496 39238
rect 21272 38344 21324 38350
rect 21272 38286 21324 38292
rect 21456 38344 21508 38350
rect 21456 38286 21508 38292
rect 21180 31748 21232 31754
rect 21180 31690 21232 31696
rect 21192 31482 21220 31690
rect 21180 31476 21232 31482
rect 21180 31418 21232 31424
rect 21180 29504 21232 29510
rect 21180 29446 21232 29452
rect 21192 28558 21220 29446
rect 21180 28552 21232 28558
rect 21180 28494 21232 28500
rect 21180 28416 21232 28422
rect 21180 28358 21232 28364
rect 21284 28370 21312 38286
rect 21364 36576 21416 36582
rect 21364 36518 21416 36524
rect 21376 36174 21404 36518
rect 21364 36168 21416 36174
rect 21364 36110 21416 36116
rect 21364 36032 21416 36038
rect 21364 35974 21416 35980
rect 21376 31754 21404 35974
rect 21456 35692 21508 35698
rect 21456 35634 21508 35640
rect 21468 34678 21496 35634
rect 21456 34672 21508 34678
rect 21456 34614 21508 34620
rect 21468 33402 21496 34614
rect 21560 33590 21588 40054
rect 21640 35556 21692 35562
rect 21640 35498 21692 35504
rect 21652 35222 21680 35498
rect 21744 35290 21772 44746
rect 22652 43988 22704 43994
rect 22652 43930 22704 43936
rect 22008 43784 22060 43790
rect 22008 43726 22060 43732
rect 22020 42226 22048 43726
rect 22664 43722 22692 43930
rect 22652 43716 22704 43722
rect 22652 43658 22704 43664
rect 22100 43648 22152 43654
rect 22100 43590 22152 43596
rect 22112 42634 22140 43590
rect 22100 42628 22152 42634
rect 22100 42570 22152 42576
rect 22652 42628 22704 42634
rect 22652 42570 22704 42576
rect 22008 42220 22060 42226
rect 22008 42162 22060 42168
rect 22020 41818 22048 42162
rect 22008 41812 22060 41818
rect 22008 41754 22060 41760
rect 22020 41414 22048 41754
rect 21928 41386 22048 41414
rect 22112 41414 22140 42570
rect 22664 42022 22692 42570
rect 22836 42560 22888 42566
rect 22836 42502 22888 42508
rect 22652 42016 22704 42022
rect 22652 41958 22704 41964
rect 22112 41386 22416 41414
rect 21824 41200 21876 41206
rect 21824 41142 21876 41148
rect 21836 40458 21864 41142
rect 21928 41070 21956 41386
rect 22284 41200 22336 41206
rect 22006 41168 22062 41177
rect 22006 41103 22008 41112
rect 22060 41103 22062 41112
rect 22282 41168 22284 41177
rect 22336 41168 22338 41177
rect 22282 41103 22338 41112
rect 22008 41074 22060 41080
rect 21916 41064 21968 41070
rect 21916 41006 21968 41012
rect 21824 40452 21876 40458
rect 21824 40394 21876 40400
rect 21928 39438 21956 41006
rect 22008 40520 22060 40526
rect 22008 40462 22060 40468
rect 22284 40520 22336 40526
rect 22284 40462 22336 40468
rect 21916 39432 21968 39438
rect 21916 39374 21968 39380
rect 21928 39030 21956 39374
rect 21916 39024 21968 39030
rect 21916 38966 21968 38972
rect 22020 38536 22048 40462
rect 22296 40050 22324 40462
rect 22284 40044 22336 40050
rect 22284 39986 22336 39992
rect 22192 39364 22244 39370
rect 22192 39306 22244 39312
rect 22100 39296 22152 39302
rect 22100 39238 22152 39244
rect 21928 38508 22048 38536
rect 21928 38350 21956 38508
rect 22006 38448 22062 38457
rect 22006 38383 22008 38392
rect 22060 38383 22062 38392
rect 22008 38354 22060 38360
rect 21824 38344 21876 38350
rect 21824 38286 21876 38292
rect 21916 38344 21968 38350
rect 21916 38286 21968 38292
rect 21836 37670 21864 38286
rect 22008 38208 22060 38214
rect 22008 38150 22060 38156
rect 22020 37874 22048 38150
rect 22112 37942 22140 39238
rect 22204 38486 22232 39306
rect 22284 39024 22336 39030
rect 22284 38966 22336 38972
rect 22296 38554 22324 38966
rect 22284 38548 22336 38554
rect 22284 38490 22336 38496
rect 22192 38480 22244 38486
rect 22192 38422 22244 38428
rect 22100 37936 22152 37942
rect 22100 37878 22152 37884
rect 22008 37868 22060 37874
rect 22008 37810 22060 37816
rect 21824 37664 21876 37670
rect 21824 37606 21876 37612
rect 21732 35284 21784 35290
rect 21732 35226 21784 35232
rect 21640 35216 21692 35222
rect 21836 35170 21864 37606
rect 21916 35760 21968 35766
rect 21916 35702 21968 35708
rect 21928 35290 21956 35702
rect 21916 35284 21968 35290
rect 21916 35226 21968 35232
rect 21640 35158 21692 35164
rect 21652 34746 21680 35158
rect 21744 35142 21864 35170
rect 21640 34740 21692 34746
rect 21640 34682 21692 34688
rect 21640 33992 21692 33998
rect 21640 33934 21692 33940
rect 21652 33658 21680 33934
rect 21640 33652 21692 33658
rect 21640 33594 21692 33600
rect 21548 33584 21600 33590
rect 21548 33526 21600 33532
rect 21744 33436 21772 35142
rect 21824 34672 21876 34678
rect 21824 34614 21876 34620
rect 21836 34542 21864 34614
rect 21824 34536 21876 34542
rect 21824 34478 21876 34484
rect 21836 34082 21864 34478
rect 21836 34054 21956 34082
rect 21824 33992 21876 33998
rect 21824 33934 21876 33940
rect 21836 33590 21864 33934
rect 21824 33584 21876 33590
rect 21824 33526 21876 33532
rect 21928 33504 21956 34054
rect 22020 33998 22048 37810
rect 22112 37194 22140 37878
rect 22192 37256 22244 37262
rect 22192 37198 22244 37204
rect 22100 37188 22152 37194
rect 22100 37130 22152 37136
rect 22204 36786 22232 37198
rect 22388 36922 22416 41386
rect 22468 38480 22520 38486
rect 22468 38422 22520 38428
rect 22376 36916 22428 36922
rect 22376 36858 22428 36864
rect 22192 36780 22244 36786
rect 22192 36722 22244 36728
rect 22100 36236 22152 36242
rect 22100 36178 22152 36184
rect 22112 34746 22140 36178
rect 22480 36122 22508 38422
rect 22560 38344 22612 38350
rect 22560 38286 22612 38292
rect 22572 38010 22600 38286
rect 22560 38004 22612 38010
rect 22560 37946 22612 37952
rect 22664 36666 22692 41958
rect 22848 40390 22876 42502
rect 22836 40384 22888 40390
rect 22836 40326 22888 40332
rect 22836 38276 22888 38282
rect 22836 38218 22888 38224
rect 22848 37942 22876 38218
rect 22836 37936 22888 37942
rect 22836 37878 22888 37884
rect 22572 36638 22692 36666
rect 22572 36310 22600 36638
rect 22940 36530 22968 45222
rect 23020 44872 23072 44878
rect 23020 44814 23072 44820
rect 22664 36502 22968 36530
rect 22560 36304 22612 36310
rect 22560 36246 22612 36252
rect 22388 36094 22508 36122
rect 22560 36100 22612 36106
rect 22192 36032 22244 36038
rect 22192 35974 22244 35980
rect 22204 35154 22232 35974
rect 22192 35148 22244 35154
rect 22192 35090 22244 35096
rect 22388 34898 22416 36094
rect 22560 36042 22612 36048
rect 22468 36032 22520 36038
rect 22468 35974 22520 35980
rect 22480 35630 22508 35974
rect 22468 35624 22520 35630
rect 22468 35566 22520 35572
rect 22468 35488 22520 35494
rect 22468 35430 22520 35436
rect 22480 35086 22508 35430
rect 22468 35080 22520 35086
rect 22468 35022 22520 35028
rect 22572 35018 22600 36042
rect 22560 35012 22612 35018
rect 22560 34954 22612 34960
rect 22388 34870 22600 34898
rect 22100 34740 22152 34746
rect 22100 34682 22152 34688
rect 22100 34604 22152 34610
rect 22100 34546 22152 34552
rect 22112 34474 22140 34546
rect 22100 34468 22152 34474
rect 22100 34410 22152 34416
rect 22008 33992 22060 33998
rect 22008 33934 22060 33940
rect 22468 33856 22520 33862
rect 22468 33798 22520 33804
rect 22284 33516 22336 33522
rect 21928 33476 22048 33504
rect 21744 33408 21864 33436
rect 21468 33374 21588 33402
rect 21376 31726 21496 31754
rect 21192 25401 21220 28358
rect 21284 28342 21404 28370
rect 21376 27577 21404 28342
rect 21362 27568 21418 27577
rect 21362 27503 21418 27512
rect 21272 27464 21324 27470
rect 21272 27406 21324 27412
rect 21364 27464 21416 27470
rect 21364 27406 21416 27412
rect 21284 26994 21312 27406
rect 21272 26988 21324 26994
rect 21272 26930 21324 26936
rect 21284 26042 21312 26930
rect 21272 26036 21324 26042
rect 21272 25978 21324 25984
rect 21178 25392 21234 25401
rect 21178 25327 21234 25336
rect 21192 24954 21220 25327
rect 21180 24948 21232 24954
rect 21180 24890 21232 24896
rect 21180 24132 21232 24138
rect 21180 24074 21232 24080
rect 21192 23322 21220 24074
rect 21180 23316 21232 23322
rect 21180 23258 21232 23264
rect 21180 22976 21232 22982
rect 21180 22918 21232 22924
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 20824 19094 21036 19122
rect 20824 18465 20852 19094
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 20810 18456 20866 18465
rect 20810 18391 20866 18400
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20718 18184 20774 18193
rect 20718 18119 20774 18128
rect 20718 18048 20774 18057
rect 20718 17983 20774 17992
rect 20732 17882 20760 17983
rect 20824 17921 20852 18226
rect 20916 18154 20944 18906
rect 21192 18714 21220 22918
rect 21272 21072 21324 21078
rect 21272 21014 21324 21020
rect 21100 18686 21220 18714
rect 21100 18408 21128 18686
rect 21180 18624 21232 18630
rect 21180 18566 21232 18572
rect 21008 18380 21128 18408
rect 20904 18148 20956 18154
rect 20904 18090 20956 18096
rect 20810 17912 20866 17921
rect 20720 17876 20772 17882
rect 20810 17847 20866 17856
rect 20720 17818 20772 17824
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20732 17241 20760 17614
rect 20824 17338 20852 17847
rect 20812 17332 20864 17338
rect 20812 17274 20864 17280
rect 20718 17232 20774 17241
rect 20718 17167 20774 17176
rect 20720 17128 20772 17134
rect 20916 17116 20944 18090
rect 20772 17088 20944 17116
rect 20720 17070 20772 17076
rect 20536 16584 20588 16590
rect 20536 16526 20588 16532
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20640 15706 20668 16050
rect 20628 15700 20680 15706
rect 20628 15642 20680 15648
rect 20444 15564 20496 15570
rect 20444 15506 20496 15512
rect 20442 15464 20498 15473
rect 20442 15399 20498 15408
rect 20456 14618 20484 15399
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20444 14612 20496 14618
rect 20444 14554 20496 14560
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20456 14074 20484 14350
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 20364 13926 20484 13954
rect 20352 13864 20404 13870
rect 20352 13806 20404 13812
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20272 11014 20300 11290
rect 20260 11008 20312 11014
rect 20260 10950 20312 10956
rect 20088 10662 20208 10690
rect 19984 10464 20036 10470
rect 19984 10406 20036 10412
rect 19340 10056 19392 10062
rect 19260 10004 19340 10010
rect 19260 9998 19392 10004
rect 19260 9982 19380 9998
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 19168 8090 19196 9522
rect 19260 8974 19288 9982
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19352 8974 19380 9318
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19156 8084 19208 8090
rect 19156 8026 19208 8032
rect 19156 7948 19208 7954
rect 19156 7890 19208 7896
rect 18892 4406 19104 4434
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18340 2746 18460 2774
rect 18236 2440 18288 2446
rect 18236 2382 18288 2388
rect 18144 2372 18196 2378
rect 18144 2314 18196 2320
rect 18340 800 18368 2746
rect 18892 2582 18920 4406
rect 19168 4282 19196 7890
rect 19260 5778 19288 8910
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 19628 7954 19656 8434
rect 19616 7948 19668 7954
rect 19616 7890 19668 7896
rect 19432 7812 19484 7818
rect 19432 7754 19484 7760
rect 19444 7274 19472 7754
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19432 7268 19484 7274
rect 19432 7210 19484 7216
rect 19444 7002 19472 7210
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19536 6798 19564 7142
rect 19524 6792 19576 6798
rect 19522 6760 19524 6769
rect 19576 6760 19578 6769
rect 19522 6695 19578 6704
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 19248 5772 19300 5778
rect 19248 5714 19300 5720
rect 19340 5636 19392 5642
rect 19340 5578 19392 5584
rect 19248 5228 19300 5234
rect 19248 5170 19300 5176
rect 19260 4622 19288 5170
rect 19352 4826 19380 5578
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 19156 4276 19208 4282
rect 19156 4218 19208 4224
rect 19444 4196 19472 5850
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19996 5166 20024 5510
rect 20088 5370 20116 10662
rect 20364 9674 20392 13806
rect 20168 9648 20220 9654
rect 20168 9590 20220 9596
rect 20272 9646 20392 9674
rect 20180 8430 20208 9590
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 20272 6644 20300 9646
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 20364 6730 20392 7142
rect 20352 6724 20404 6730
rect 20352 6666 20404 6672
rect 20263 6616 20300 6644
rect 20263 6474 20291 6616
rect 20168 6452 20220 6458
rect 20263 6446 20300 6474
rect 20168 6394 20220 6400
rect 20180 5914 20208 6394
rect 20168 5908 20220 5914
rect 20168 5850 20220 5856
rect 20076 5364 20128 5370
rect 20076 5306 20128 5312
rect 20168 5296 20220 5302
rect 20168 5238 20220 5244
rect 19984 5160 20036 5166
rect 19984 5102 20036 5108
rect 19708 5092 19760 5098
rect 19708 5034 19760 5040
rect 19720 4729 19748 5034
rect 19706 4720 19762 4729
rect 19706 4655 19762 4664
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19352 4168 19472 4196
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19156 4072 19208 4078
rect 19156 4014 19208 4020
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 18880 2576 18932 2582
rect 18880 2518 18932 2524
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 18708 800 18736 2246
rect 19076 800 19104 3538
rect 19168 3194 19196 4014
rect 19260 3738 19288 4082
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 19248 3392 19300 3398
rect 19248 3334 19300 3340
rect 19156 3188 19208 3194
rect 19156 3130 19208 3136
rect 19260 2990 19288 3334
rect 19248 2984 19300 2990
rect 19248 2926 19300 2932
rect 19352 1442 19380 4168
rect 19616 4004 19668 4010
rect 19616 3946 19668 3952
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19444 3176 19472 3470
rect 19536 3466 19564 3878
rect 19628 3602 19656 3946
rect 19892 3664 19944 3670
rect 19892 3606 19944 3612
rect 19616 3596 19668 3602
rect 19616 3538 19668 3544
rect 19904 3505 19932 3606
rect 19890 3496 19946 3505
rect 19524 3460 19576 3466
rect 19890 3431 19946 3440
rect 19524 3402 19576 3408
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19444 3148 19564 3176
rect 19432 2848 19484 2854
rect 19432 2790 19484 2796
rect 19444 2446 19472 2790
rect 19536 2650 19564 3148
rect 19996 3126 20024 4422
rect 20088 4010 20116 4558
rect 20076 4004 20128 4010
rect 20076 3946 20128 3952
rect 19984 3120 20036 3126
rect 19984 3062 20036 3068
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 20076 2304 20128 2310
rect 20076 2246 20128 2252
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19352 1414 19472 1442
rect 19444 800 19472 1414
rect 19812 870 19932 898
rect 19812 800 19840 870
rect 202 0 258 800
rect 570 0 626 800
rect 938 0 994 800
rect 1306 0 1362 800
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13542 0 13598 800
rect 13910 0 13966 800
rect 14278 0 14334 800
rect 14646 0 14702 800
rect 15014 0 15070 800
rect 15382 0 15438 800
rect 15750 0 15806 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16854 0 16910 800
rect 17222 0 17278 800
rect 17590 0 17646 800
rect 17958 0 18014 800
rect 18326 0 18382 800
rect 18694 0 18750 800
rect 19062 0 19118 800
rect 19430 0 19486 800
rect 19798 0 19854 800
rect 19904 762 19932 870
rect 20088 762 20116 2246
rect 20180 800 20208 5238
rect 20272 2378 20300 6446
rect 20352 5568 20404 5574
rect 20352 5510 20404 5516
rect 20364 4078 20392 5510
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 20352 3936 20404 3942
rect 20352 3878 20404 3884
rect 20364 2990 20392 3878
rect 20352 2984 20404 2990
rect 20352 2926 20404 2932
rect 20456 2378 20484 13926
rect 20548 13394 20576 14894
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20548 11830 20576 12786
rect 20732 12730 20760 15302
rect 20640 12702 20760 12730
rect 20640 12209 20668 12702
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20626 12200 20682 12209
rect 20732 12170 20760 12582
rect 20626 12135 20682 12144
rect 20720 12164 20772 12170
rect 20720 12106 20772 12112
rect 20824 12050 20852 16526
rect 21008 16130 21036 18380
rect 21086 18320 21142 18329
rect 21086 18255 21142 18264
rect 20916 16102 21036 16130
rect 20916 15978 20944 16102
rect 21100 15994 21128 18255
rect 20904 15972 20956 15978
rect 20904 15914 20956 15920
rect 21008 15966 21128 15994
rect 21008 15162 21036 15966
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 21100 15502 21128 15846
rect 21088 15496 21140 15502
rect 21088 15438 21140 15444
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 20904 14612 20956 14618
rect 20904 14554 20956 14560
rect 20916 14278 20944 14554
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 20916 12714 20944 14214
rect 20904 12708 20956 12714
rect 20904 12650 20956 12656
rect 20640 12022 20852 12050
rect 20536 11824 20588 11830
rect 20536 11766 20588 11772
rect 20536 11076 20588 11082
rect 20536 11018 20588 11024
rect 20548 8634 20576 11018
rect 20640 9654 20668 12022
rect 21088 11756 21140 11762
rect 21088 11698 21140 11704
rect 21100 11354 21128 11698
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 21088 11144 21140 11150
rect 21088 11086 21140 11092
rect 21100 10810 21128 11086
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 20904 9988 20956 9994
rect 20904 9930 20956 9936
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20628 9648 20680 9654
rect 20628 9590 20680 9596
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 20732 7886 20760 9862
rect 20916 9722 20944 9930
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20536 7404 20588 7410
rect 20536 7346 20588 7352
rect 20548 6458 20576 7346
rect 21086 6760 21142 6769
rect 21086 6695 21142 6704
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20640 6458 20668 6598
rect 20536 6452 20588 6458
rect 20536 6394 20588 6400
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 21100 6322 21128 6695
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 21100 5846 21128 6258
rect 21088 5840 21140 5846
rect 21088 5782 21140 5788
rect 20536 5636 20588 5642
rect 20536 5578 20588 5584
rect 20260 2372 20312 2378
rect 20260 2314 20312 2320
rect 20444 2372 20496 2378
rect 20444 2314 20496 2320
rect 20548 800 20576 5578
rect 20996 5092 21048 5098
rect 20996 5034 21048 5040
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20810 4856 20866 4865
rect 20810 4791 20866 4800
rect 20824 4758 20852 4791
rect 20812 4752 20864 4758
rect 20812 4694 20864 4700
rect 20916 4690 20944 4966
rect 20904 4684 20956 4690
rect 20904 4626 20956 4632
rect 20904 3936 20956 3942
rect 20904 3878 20956 3884
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20732 3058 20760 3674
rect 20916 3466 20944 3878
rect 20904 3460 20956 3466
rect 20904 3402 20956 3408
rect 21008 3058 21036 5034
rect 21100 4282 21128 5782
rect 21088 4276 21140 4282
rect 21088 4218 21140 4224
rect 21088 4140 21140 4146
rect 21088 4082 21140 4088
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20996 3052 21048 3058
rect 20996 2994 21048 3000
rect 20812 2848 20864 2854
rect 20812 2790 20864 2796
rect 20824 2446 20852 2790
rect 21100 2650 21128 4082
rect 21088 2644 21140 2650
rect 21088 2586 21140 2592
rect 20904 2576 20956 2582
rect 20904 2518 20956 2524
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 20916 800 20944 2518
rect 21192 2378 21220 18566
rect 21284 18329 21312 21014
rect 21376 20505 21404 27406
rect 21362 20496 21418 20505
rect 21362 20431 21418 20440
rect 21270 18320 21326 18329
rect 21270 18255 21326 18264
rect 21272 18148 21324 18154
rect 21272 18090 21324 18096
rect 21284 17610 21312 18090
rect 21272 17604 21324 17610
rect 21272 17546 21324 17552
rect 21272 15496 21324 15502
rect 21272 15438 21324 15444
rect 21284 15162 21312 15438
rect 21272 15156 21324 15162
rect 21272 15098 21324 15104
rect 21284 15026 21312 15098
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 21272 12844 21324 12850
rect 21272 12786 21324 12792
rect 21284 11762 21312 12786
rect 21376 11898 21404 20431
rect 21468 18766 21496 31726
rect 21560 29034 21588 33374
rect 21836 31754 21864 33408
rect 22020 31958 22048 33476
rect 22284 33458 22336 33464
rect 22192 33448 22244 33454
rect 22192 33390 22244 33396
rect 22100 32904 22152 32910
rect 22100 32846 22152 32852
rect 22112 32570 22140 32846
rect 22100 32564 22152 32570
rect 22100 32506 22152 32512
rect 22100 32360 22152 32366
rect 22100 32302 22152 32308
rect 22008 31952 22060 31958
rect 22008 31894 22060 31900
rect 21732 31748 21784 31754
rect 21836 31726 21956 31754
rect 21732 31690 21784 31696
rect 21640 30388 21692 30394
rect 21640 30330 21692 30336
rect 21548 29028 21600 29034
rect 21548 28970 21600 28976
rect 21548 28688 21600 28694
rect 21548 28630 21600 28636
rect 21560 28558 21588 28630
rect 21548 28552 21600 28558
rect 21548 28494 21600 28500
rect 21560 28014 21588 28494
rect 21548 28008 21600 28014
rect 21548 27950 21600 27956
rect 21548 25900 21600 25906
rect 21548 25842 21600 25848
rect 21560 25294 21588 25842
rect 21652 25838 21680 30330
rect 21744 27316 21772 31690
rect 21824 31476 21876 31482
rect 21824 31418 21876 31424
rect 21836 30326 21864 31418
rect 21824 30320 21876 30326
rect 21824 30262 21876 30268
rect 21928 29322 21956 31726
rect 22020 31278 22048 31894
rect 22112 31754 22140 32302
rect 22204 31890 22232 33390
rect 22296 33114 22324 33458
rect 22284 33108 22336 33114
rect 22284 33050 22336 33056
rect 22192 31884 22244 31890
rect 22192 31826 22244 31832
rect 22100 31748 22152 31754
rect 22100 31690 22152 31696
rect 22100 31340 22152 31346
rect 22100 31282 22152 31288
rect 22008 31272 22060 31278
rect 22008 31214 22060 31220
rect 22112 30394 22140 31282
rect 22100 30388 22152 30394
rect 22100 30330 22152 30336
rect 22204 30190 22232 31826
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 22296 30734 22324 31282
rect 22284 30728 22336 30734
rect 22284 30670 22336 30676
rect 22284 30592 22336 30598
rect 22284 30534 22336 30540
rect 22192 30184 22244 30190
rect 22192 30126 22244 30132
rect 22204 29850 22232 30126
rect 22192 29844 22244 29850
rect 22192 29786 22244 29792
rect 21836 29294 21956 29322
rect 22008 29300 22060 29306
rect 21836 28529 21864 29294
rect 22008 29242 22060 29248
rect 21916 29232 21968 29238
rect 21916 29174 21968 29180
rect 21822 28520 21878 28529
rect 21822 28455 21878 28464
rect 21824 28416 21876 28422
rect 21824 28358 21876 28364
rect 21836 27470 21864 28358
rect 21928 28082 21956 29174
rect 22020 28694 22048 29242
rect 22204 29238 22232 29786
rect 22192 29232 22244 29238
rect 22192 29174 22244 29180
rect 22100 29164 22152 29170
rect 22100 29106 22152 29112
rect 22112 28762 22140 29106
rect 22100 28756 22152 28762
rect 22100 28698 22152 28704
rect 22008 28688 22060 28694
rect 22008 28630 22060 28636
rect 22006 28520 22062 28529
rect 22006 28455 22062 28464
rect 21916 28076 21968 28082
rect 21916 28018 21968 28024
rect 21824 27464 21876 27470
rect 21824 27406 21876 27412
rect 21744 27288 21864 27316
rect 21732 26920 21784 26926
rect 21732 26862 21784 26868
rect 21744 26518 21772 26862
rect 21732 26512 21784 26518
rect 21732 26454 21784 26460
rect 21640 25832 21692 25838
rect 21640 25774 21692 25780
rect 21548 25288 21600 25294
rect 21548 25230 21600 25236
rect 21560 24206 21588 25230
rect 21548 24200 21600 24206
rect 21548 24142 21600 24148
rect 21652 24138 21680 25774
rect 21640 24132 21692 24138
rect 21640 24074 21692 24080
rect 21548 22228 21600 22234
rect 21548 22170 21600 22176
rect 21447 18760 21499 18766
rect 21447 18702 21499 18708
rect 21468 18222 21496 18702
rect 21456 18216 21508 18222
rect 21456 18158 21508 18164
rect 21456 17196 21508 17202
rect 21456 17138 21508 17144
rect 21468 16726 21496 17138
rect 21456 16720 21508 16726
rect 21456 16662 21508 16668
rect 21560 13938 21588 22170
rect 21732 21888 21784 21894
rect 21732 21830 21784 21836
rect 21744 20330 21772 21830
rect 21732 20324 21784 20330
rect 21732 20266 21784 20272
rect 21744 19922 21772 20266
rect 21732 19916 21784 19922
rect 21732 19858 21784 19864
rect 21640 18896 21692 18902
rect 21640 18838 21692 18844
rect 21652 18290 21680 18838
rect 21640 18284 21692 18290
rect 21640 18226 21692 18232
rect 21732 18080 21784 18086
rect 21732 18022 21784 18028
rect 21744 17678 21772 18022
rect 21732 17672 21784 17678
rect 21732 17614 21784 17620
rect 21640 17536 21692 17542
rect 21640 17478 21692 17484
rect 21652 17134 21680 17478
rect 21640 17128 21692 17134
rect 21640 17070 21692 17076
rect 21652 16590 21680 17070
rect 21640 16584 21692 16590
rect 21640 16526 21692 16532
rect 21732 16584 21784 16590
rect 21732 16526 21784 16532
rect 21744 16250 21772 16526
rect 21732 16244 21784 16250
rect 21732 16186 21784 16192
rect 21548 13932 21600 13938
rect 21548 13874 21600 13880
rect 21560 13462 21588 13874
rect 21548 13456 21600 13462
rect 21548 13398 21600 13404
rect 21836 12434 21864 27288
rect 22020 25498 22048 28455
rect 22296 28200 22324 30534
rect 22480 30376 22508 33798
rect 22112 28172 22324 28200
rect 22388 30348 22508 30376
rect 22008 25492 22060 25498
rect 22008 25434 22060 25440
rect 22112 24954 22140 28172
rect 22192 28076 22244 28082
rect 22192 28018 22244 28024
rect 22204 27606 22232 28018
rect 22192 27600 22244 27606
rect 22192 27542 22244 27548
rect 22284 27464 22336 27470
rect 22204 27424 22284 27452
rect 22100 24948 22152 24954
rect 22100 24890 22152 24896
rect 22100 24200 22152 24206
rect 22100 24142 22152 24148
rect 22006 23896 22062 23905
rect 22006 23831 22062 23840
rect 22020 23526 22048 23831
rect 22112 23730 22140 24142
rect 22100 23724 22152 23730
rect 22100 23666 22152 23672
rect 22100 23588 22152 23594
rect 22100 23530 22152 23536
rect 22008 23520 22060 23526
rect 22008 23462 22060 23468
rect 21916 22976 21968 22982
rect 21916 22918 21968 22924
rect 21928 22642 21956 22918
rect 21916 22636 21968 22642
rect 21916 22578 21968 22584
rect 22112 22094 22140 23530
rect 22204 23254 22232 27424
rect 22284 27406 22336 27412
rect 22284 27328 22336 27334
rect 22284 27270 22336 27276
rect 22296 26994 22324 27270
rect 22284 26988 22336 26994
rect 22284 26930 22336 26936
rect 22284 26852 22336 26858
rect 22284 26794 22336 26800
rect 22296 23594 22324 26794
rect 22284 23588 22336 23594
rect 22284 23530 22336 23536
rect 22192 23248 22244 23254
rect 22192 23190 22244 23196
rect 22204 22982 22232 23190
rect 22284 23112 22336 23118
rect 22284 23054 22336 23060
rect 22192 22976 22244 22982
rect 22192 22918 22244 22924
rect 22112 22066 22232 22094
rect 22100 21956 22152 21962
rect 22100 21898 22152 21904
rect 22112 21350 22140 21898
rect 22100 21344 22152 21350
rect 22100 21286 22152 21292
rect 22008 20460 22060 20466
rect 22008 20402 22060 20408
rect 22020 19922 22048 20402
rect 22008 19916 22060 19922
rect 22008 19858 22060 19864
rect 22020 19334 22048 19858
rect 21928 19306 22048 19334
rect 21928 18290 21956 19306
rect 22112 18902 22140 21286
rect 22204 20074 22232 22066
rect 22296 21146 22324 23054
rect 22388 21978 22416 30348
rect 22468 29640 22520 29646
rect 22468 29582 22520 29588
rect 22480 29170 22508 29582
rect 22468 29164 22520 29170
rect 22468 29106 22520 29112
rect 22468 28960 22520 28966
rect 22468 28902 22520 28908
rect 22480 28558 22508 28902
rect 22468 28552 22520 28558
rect 22468 28494 22520 28500
rect 22468 25288 22520 25294
rect 22468 25230 22520 25236
rect 22480 22710 22508 25230
rect 22572 24886 22600 34870
rect 22664 28665 22692 36502
rect 22928 36100 22980 36106
rect 22928 36042 22980 36048
rect 22744 35760 22796 35766
rect 22744 35702 22796 35708
rect 22756 34746 22784 35702
rect 22940 35698 22968 36042
rect 22928 35692 22980 35698
rect 22928 35634 22980 35640
rect 22744 34740 22796 34746
rect 22744 34682 22796 34688
rect 22836 34468 22888 34474
rect 22836 34410 22888 34416
rect 22744 32904 22796 32910
rect 22742 32872 22744 32881
rect 22796 32872 22798 32881
rect 22742 32807 22798 32816
rect 22744 32564 22796 32570
rect 22744 32506 22796 32512
rect 22756 30598 22784 32506
rect 22744 30592 22796 30598
rect 22744 30534 22796 30540
rect 22744 29776 22796 29782
rect 22744 29718 22796 29724
rect 22756 29578 22784 29718
rect 22744 29572 22796 29578
rect 22744 29514 22796 29520
rect 22848 29306 22876 34410
rect 22928 30796 22980 30802
rect 22928 30738 22980 30744
rect 22836 29300 22888 29306
rect 22836 29242 22888 29248
rect 22650 28656 22706 28665
rect 22940 28642 22968 30738
rect 22650 28591 22706 28600
rect 22848 28614 22968 28642
rect 22848 26994 22876 28614
rect 22928 28484 22980 28490
rect 22928 28426 22980 28432
rect 22940 28121 22968 28426
rect 22926 28112 22982 28121
rect 22926 28047 22982 28056
rect 23032 27470 23060 44814
rect 23296 43784 23348 43790
rect 23296 43726 23348 43732
rect 23308 42650 23336 43726
rect 23400 42770 23428 46922
rect 23480 44328 23532 44334
rect 23480 44270 23532 44276
rect 23388 42764 23440 42770
rect 23388 42706 23440 42712
rect 23308 42622 23428 42650
rect 23204 40180 23256 40186
rect 23204 40122 23256 40128
rect 23216 39982 23244 40122
rect 23204 39976 23256 39982
rect 23204 39918 23256 39924
rect 23216 38554 23244 39918
rect 23296 39908 23348 39914
rect 23296 39850 23348 39856
rect 23204 38548 23256 38554
rect 23204 38490 23256 38496
rect 23112 38344 23164 38350
rect 23164 38304 23244 38332
rect 23112 38286 23164 38292
rect 23112 31748 23164 31754
rect 23112 31690 23164 31696
rect 23124 30938 23152 31690
rect 23112 30932 23164 30938
rect 23112 30874 23164 30880
rect 23112 30252 23164 30258
rect 23112 30194 23164 30200
rect 23124 29850 23152 30194
rect 23112 29844 23164 29850
rect 23112 29786 23164 29792
rect 23216 27690 23244 38304
rect 23308 37398 23336 39850
rect 23400 37398 23428 42622
rect 23492 39914 23520 44270
rect 23952 43450 23980 46922
rect 24032 46572 24084 46578
rect 24032 46514 24084 46520
rect 24044 45558 24072 46514
rect 24032 45552 24084 45558
rect 24032 45494 24084 45500
rect 24216 45484 24268 45490
rect 24216 45426 24268 45432
rect 24032 44396 24084 44402
rect 24032 44338 24084 44344
rect 24044 43994 24072 44338
rect 24032 43988 24084 43994
rect 24032 43930 24084 43936
rect 23940 43444 23992 43450
rect 23940 43386 23992 43392
rect 24124 43308 24176 43314
rect 24124 43250 24176 43256
rect 24136 42362 24164 43250
rect 24124 42356 24176 42362
rect 24124 42298 24176 42304
rect 24032 42220 24084 42226
rect 24032 42162 24084 42168
rect 23848 42152 23900 42158
rect 23848 42094 23900 42100
rect 23860 41002 23888 42094
rect 24044 41750 24072 42162
rect 24032 41744 24084 41750
rect 24032 41686 24084 41692
rect 23848 40996 23900 41002
rect 23848 40938 23900 40944
rect 23480 39908 23532 39914
rect 23480 39850 23532 39856
rect 23756 38752 23808 38758
rect 23756 38694 23808 38700
rect 23768 38350 23796 38694
rect 23756 38344 23808 38350
rect 23756 38286 23808 38292
rect 23296 37392 23348 37398
rect 23296 37334 23348 37340
rect 23388 37392 23440 37398
rect 23388 37334 23440 37340
rect 23308 36922 23336 37334
rect 23756 37120 23808 37126
rect 23756 37062 23808 37068
rect 23768 36922 23796 37062
rect 23296 36916 23348 36922
rect 23296 36858 23348 36864
rect 23756 36916 23808 36922
rect 23756 36858 23808 36864
rect 23388 36780 23440 36786
rect 23388 36722 23440 36728
rect 23664 36780 23716 36786
rect 23664 36722 23716 36728
rect 23296 34468 23348 34474
rect 23296 34410 23348 34416
rect 23308 33998 23336 34410
rect 23296 33992 23348 33998
rect 23296 33934 23348 33940
rect 23308 33658 23336 33934
rect 23296 33652 23348 33658
rect 23296 33594 23348 33600
rect 23296 32836 23348 32842
rect 23296 32778 23348 32784
rect 23308 32570 23336 32778
rect 23296 32564 23348 32570
rect 23296 32506 23348 32512
rect 23296 31136 23348 31142
rect 23296 31078 23348 31084
rect 23308 30734 23336 31078
rect 23296 30728 23348 30734
rect 23296 30670 23348 30676
rect 23296 29640 23348 29646
rect 23294 29608 23296 29617
rect 23348 29608 23350 29617
rect 23294 29543 23350 29552
rect 23296 29028 23348 29034
rect 23296 28970 23348 28976
rect 23308 28762 23336 28970
rect 23296 28756 23348 28762
rect 23296 28698 23348 28704
rect 23296 28484 23348 28490
rect 23296 28426 23348 28432
rect 23124 27662 23244 27690
rect 23020 27464 23072 27470
rect 23020 27406 23072 27412
rect 22836 26988 22888 26994
rect 22836 26930 22888 26936
rect 23124 26874 23152 27662
rect 23308 27606 23336 28426
rect 23400 27946 23428 36722
rect 23676 36650 23704 36722
rect 23664 36644 23716 36650
rect 23664 36586 23716 36592
rect 23572 34944 23624 34950
rect 23572 34886 23624 34892
rect 23584 34678 23612 34886
rect 23572 34672 23624 34678
rect 23572 34614 23624 34620
rect 23676 34082 23704 36586
rect 23940 35012 23992 35018
rect 23940 34954 23992 34960
rect 23848 34944 23900 34950
rect 23848 34886 23900 34892
rect 23860 34202 23888 34886
rect 23952 34542 23980 34954
rect 24228 34746 24256 45426
rect 24412 44538 24440 46990
rect 24504 46918 24532 49200
rect 25332 47258 25360 49200
rect 25320 47252 25372 47258
rect 25320 47194 25372 47200
rect 24584 46980 24636 46986
rect 24584 46922 24636 46928
rect 24492 46912 24544 46918
rect 24492 46854 24544 46860
rect 24400 44532 24452 44538
rect 24400 44474 24452 44480
rect 24596 43450 24624 46922
rect 26160 46714 26188 49200
rect 27080 47054 27108 49200
rect 27528 47660 27580 47666
rect 27528 47602 27580 47608
rect 27540 47258 27568 47602
rect 27528 47252 27580 47258
rect 27528 47194 27580 47200
rect 27068 47048 27120 47054
rect 27068 46990 27120 46996
rect 27908 46986 27936 49200
rect 28172 47116 28224 47122
rect 28920 47104 28948 49286
rect 29550 49286 29684 49314
rect 29550 49200 29606 49286
rect 29000 47116 29052 47122
rect 28920 47076 29000 47104
rect 28172 47058 28224 47064
rect 29000 47058 29052 47064
rect 27896 46980 27948 46986
rect 27896 46922 27948 46928
rect 26148 46708 26200 46714
rect 26148 46650 26200 46656
rect 25044 45008 25096 45014
rect 25044 44950 25096 44956
rect 24584 43444 24636 43450
rect 24584 43386 24636 43392
rect 24768 43308 24820 43314
rect 24768 43250 24820 43256
rect 24780 42906 24808 43250
rect 24768 42900 24820 42906
rect 24768 42842 24820 42848
rect 25056 40050 25084 44950
rect 27712 42764 27764 42770
rect 27712 42706 27764 42712
rect 27528 42220 27580 42226
rect 27528 42162 27580 42168
rect 27540 41818 27568 42162
rect 27528 41812 27580 41818
rect 27528 41754 27580 41760
rect 27252 41540 27304 41546
rect 27252 41482 27304 41488
rect 25412 40724 25464 40730
rect 25412 40666 25464 40672
rect 24860 40044 24912 40050
rect 24860 39986 24912 39992
rect 25044 40044 25096 40050
rect 25044 39986 25096 39992
rect 24308 39840 24360 39846
rect 24308 39782 24360 39788
rect 24320 37466 24348 39782
rect 24872 39642 24900 39986
rect 25424 39642 25452 40666
rect 25504 40112 25556 40118
rect 25504 40054 25556 40060
rect 24860 39636 24912 39642
rect 24860 39578 24912 39584
rect 25412 39636 25464 39642
rect 25412 39578 25464 39584
rect 25136 39568 25188 39574
rect 25136 39510 25188 39516
rect 24860 39364 24912 39370
rect 24860 39306 24912 39312
rect 24308 37460 24360 37466
rect 24308 37402 24360 37408
rect 24492 37120 24544 37126
rect 24492 37062 24544 37068
rect 24504 36786 24532 37062
rect 24492 36780 24544 36786
rect 24492 36722 24544 36728
rect 24308 36576 24360 36582
rect 24308 36518 24360 36524
rect 24320 35698 24348 36518
rect 24308 35692 24360 35698
rect 24308 35634 24360 35640
rect 24492 35488 24544 35494
rect 24492 35430 24544 35436
rect 24216 34740 24268 34746
rect 24216 34682 24268 34688
rect 23940 34536 23992 34542
rect 23940 34478 23992 34484
rect 23848 34196 23900 34202
rect 23848 34138 23900 34144
rect 23492 34054 23704 34082
rect 23492 33318 23520 34054
rect 23664 33856 23716 33862
rect 23664 33798 23716 33804
rect 23480 33312 23532 33318
rect 23480 33254 23532 33260
rect 23492 32774 23520 33254
rect 23572 32836 23624 32842
rect 23572 32778 23624 32784
rect 23480 32768 23532 32774
rect 23480 32710 23532 32716
rect 23584 32026 23612 32778
rect 23676 32570 23704 33798
rect 23664 32564 23716 32570
rect 23664 32506 23716 32512
rect 23572 32020 23624 32026
rect 23572 31962 23624 31968
rect 23664 31680 23716 31686
rect 23664 31622 23716 31628
rect 23572 31272 23624 31278
rect 23676 31260 23704 31622
rect 23624 31232 23704 31260
rect 23572 31214 23624 31220
rect 23572 30728 23624 30734
rect 23572 30670 23624 30676
rect 23584 30394 23612 30670
rect 23572 30388 23624 30394
rect 23572 30330 23624 30336
rect 23572 29640 23624 29646
rect 23572 29582 23624 29588
rect 23584 29306 23612 29582
rect 23572 29300 23624 29306
rect 23572 29242 23624 29248
rect 23480 28416 23532 28422
rect 23480 28358 23532 28364
rect 23388 27940 23440 27946
rect 23388 27882 23440 27888
rect 23296 27600 23348 27606
rect 23296 27542 23348 27548
rect 23204 27532 23256 27538
rect 23204 27474 23256 27480
rect 23216 27062 23244 27474
rect 23296 27396 23348 27402
rect 23296 27338 23348 27344
rect 23204 27056 23256 27062
rect 23204 26998 23256 27004
rect 22848 26846 23152 26874
rect 23308 26858 23336 27338
rect 23492 27334 23520 28358
rect 23570 27432 23626 27441
rect 23570 27367 23626 27376
rect 23584 27334 23612 27367
rect 23480 27328 23532 27334
rect 23480 27270 23532 27276
rect 23572 27328 23624 27334
rect 23572 27270 23624 27276
rect 23296 26852 23348 26858
rect 22744 26240 22796 26246
rect 22744 26182 22796 26188
rect 22756 25294 22784 26182
rect 22744 25288 22796 25294
rect 22744 25230 22796 25236
rect 22560 24880 22612 24886
rect 22560 24822 22612 24828
rect 22652 24812 22704 24818
rect 22652 24754 22704 24760
rect 22664 24138 22692 24754
rect 22744 24608 22796 24614
rect 22744 24550 22796 24556
rect 22652 24132 22704 24138
rect 22652 24074 22704 24080
rect 22560 23792 22612 23798
rect 22560 23734 22612 23740
rect 22572 23118 22600 23734
rect 22664 23730 22692 24074
rect 22652 23724 22704 23730
rect 22652 23666 22704 23672
rect 22560 23112 22612 23118
rect 22560 23054 22612 23060
rect 22560 22976 22612 22982
rect 22560 22918 22612 22924
rect 22468 22704 22520 22710
rect 22468 22646 22520 22652
rect 22480 22098 22508 22646
rect 22468 22092 22520 22098
rect 22468 22034 22520 22040
rect 22388 21950 22508 21978
rect 22284 21140 22336 21146
rect 22284 21082 22336 21088
rect 22204 20046 22324 20074
rect 22100 18896 22152 18902
rect 22100 18838 22152 18844
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 21916 18284 21968 18290
rect 21916 18226 21968 18232
rect 22020 18086 22048 18702
rect 22008 18080 22060 18086
rect 22008 18022 22060 18028
rect 22192 16652 22244 16658
rect 22192 16594 22244 16600
rect 22008 16244 22060 16250
rect 22008 16186 22060 16192
rect 21916 16040 21968 16046
rect 21916 15982 21968 15988
rect 21928 14618 21956 15982
rect 22020 15502 22048 16186
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 22100 15360 22152 15366
rect 22100 15302 22152 15308
rect 22112 15026 22140 15302
rect 22204 15094 22232 16594
rect 22192 15088 22244 15094
rect 22192 15030 22244 15036
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 22008 14816 22060 14822
rect 22008 14758 22060 14764
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 22020 14414 22048 14758
rect 22008 14408 22060 14414
rect 22008 14350 22060 14356
rect 22204 13938 22232 15030
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 21744 12406 21864 12434
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 21272 11756 21324 11762
rect 21272 11698 21324 11704
rect 21284 10674 21312 11698
rect 21376 11150 21404 11834
rect 21456 11620 21508 11626
rect 21456 11562 21508 11568
rect 21468 11354 21496 11562
rect 21456 11348 21508 11354
rect 21456 11290 21508 11296
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 21272 10668 21324 10674
rect 21272 10610 21324 10616
rect 21744 9926 21772 12406
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 21836 11762 21864 12174
rect 21824 11756 21876 11762
rect 21824 11698 21876 11704
rect 21916 11280 21968 11286
rect 21916 11222 21968 11228
rect 21928 10674 21956 11222
rect 21916 10668 21968 10674
rect 21916 10610 21968 10616
rect 21916 10056 21968 10062
rect 21916 9998 21968 10004
rect 21732 9920 21784 9926
rect 21732 9862 21784 9868
rect 21928 9586 21956 9998
rect 22100 9716 22152 9722
rect 22100 9658 22152 9664
rect 21548 9580 21600 9586
rect 21548 9522 21600 9528
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 21560 9178 21588 9522
rect 22112 9178 22140 9658
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 22296 9058 22324 20046
rect 22376 19712 22428 19718
rect 22376 19654 22428 19660
rect 22388 18766 22416 19654
rect 22376 18760 22428 18766
rect 22376 18702 22428 18708
rect 22480 17728 22508 21950
rect 22572 21468 22600 22918
rect 22664 21690 22692 23666
rect 22756 21865 22784 24550
rect 22848 24070 22876 26846
rect 23296 26794 23348 26800
rect 23112 26784 23164 26790
rect 23112 26726 23164 26732
rect 23124 26382 23152 26726
rect 23308 26382 23336 26794
rect 22928 26376 22980 26382
rect 22928 26318 22980 26324
rect 23112 26376 23164 26382
rect 23112 26318 23164 26324
rect 23296 26376 23348 26382
rect 23296 26318 23348 26324
rect 22836 24064 22888 24070
rect 22836 24006 22888 24012
rect 22848 23866 22876 24006
rect 22836 23860 22888 23866
rect 22836 23802 22888 23808
rect 22836 21956 22888 21962
rect 22836 21898 22888 21904
rect 22742 21856 22798 21865
rect 22742 21791 22798 21800
rect 22652 21684 22704 21690
rect 22652 21626 22704 21632
rect 22756 21622 22784 21791
rect 22848 21690 22876 21898
rect 22836 21684 22888 21690
rect 22836 21626 22888 21632
rect 22744 21616 22796 21622
rect 22744 21558 22796 21564
rect 22572 21440 22784 21468
rect 22652 20868 22704 20874
rect 22652 20810 22704 20816
rect 22664 19854 22692 20810
rect 22652 19848 22704 19854
rect 22652 19790 22704 19796
rect 22560 18284 22612 18290
rect 22560 18226 22612 18232
rect 22572 17882 22600 18226
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 22388 17700 22508 17728
rect 22388 17134 22416 17700
rect 22468 17604 22520 17610
rect 22468 17546 22520 17552
rect 22480 17338 22508 17546
rect 22560 17536 22612 17542
rect 22560 17478 22612 17484
rect 22468 17332 22520 17338
rect 22468 17274 22520 17280
rect 22376 17128 22428 17134
rect 22376 17070 22428 17076
rect 22572 16522 22600 17478
rect 22560 16516 22612 16522
rect 22560 16458 22612 16464
rect 22468 16108 22520 16114
rect 22468 16050 22520 16056
rect 22480 15978 22508 16050
rect 22468 15972 22520 15978
rect 22468 15914 22520 15920
rect 22480 15638 22508 15914
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22468 15632 22520 15638
rect 22468 15574 22520 15580
rect 22572 15570 22600 15846
rect 22560 15564 22612 15570
rect 22560 15506 22612 15512
rect 22664 9674 22692 19790
rect 22756 14414 22784 21440
rect 22744 14408 22796 14414
rect 22744 14350 22796 14356
rect 22756 14006 22784 14350
rect 22744 14000 22796 14006
rect 22744 13942 22796 13948
rect 22744 12164 22796 12170
rect 22744 12106 22796 12112
rect 22756 10742 22784 12106
rect 22744 10736 22796 10742
rect 22744 10678 22796 10684
rect 22376 9648 22428 9654
rect 22664 9646 22876 9674
rect 22376 9590 22428 9596
rect 22112 9030 22324 9058
rect 21364 8968 21416 8974
rect 21364 8910 21416 8916
rect 21270 8528 21326 8537
rect 21270 8463 21326 8472
rect 21284 8362 21312 8463
rect 21272 8356 21324 8362
rect 21272 8298 21324 8304
rect 21284 7750 21312 8298
rect 21376 8090 21404 8910
rect 21456 8900 21508 8906
rect 21456 8842 21508 8848
rect 21468 8430 21496 8842
rect 21640 8492 21692 8498
rect 21640 8434 21692 8440
rect 21732 8492 21784 8498
rect 21732 8434 21784 8440
rect 21456 8424 21508 8430
rect 21456 8366 21508 8372
rect 21468 8294 21496 8366
rect 21456 8288 21508 8294
rect 21456 8230 21508 8236
rect 21364 8084 21416 8090
rect 21364 8026 21416 8032
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 21284 7478 21312 7686
rect 21272 7472 21324 7478
rect 21272 7414 21324 7420
rect 21364 6996 21416 7002
rect 21364 6938 21416 6944
rect 21376 6390 21404 6938
rect 21364 6384 21416 6390
rect 21364 6326 21416 6332
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 21180 2372 21232 2378
rect 21180 2314 21232 2320
rect 21284 800 21312 5170
rect 21456 4072 21508 4078
rect 21456 4014 21508 4020
rect 21468 3738 21496 4014
rect 21456 3732 21508 3738
rect 21456 3674 21508 3680
rect 21652 800 21680 8434
rect 21744 7886 21772 8434
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21916 7472 21968 7478
rect 21916 7414 21968 7420
rect 21824 6656 21876 6662
rect 21824 6598 21876 6604
rect 21836 6322 21864 6598
rect 21824 6316 21876 6322
rect 21824 6258 21876 6264
rect 21928 6202 21956 7414
rect 22008 7336 22060 7342
rect 22008 7278 22060 7284
rect 22020 7002 22048 7278
rect 22008 6996 22060 7002
rect 22008 6938 22060 6944
rect 22112 6882 22140 9030
rect 22192 8900 22244 8906
rect 22192 8842 22244 8848
rect 22284 8900 22336 8906
rect 22284 8842 22336 8848
rect 22204 8537 22232 8842
rect 22190 8528 22246 8537
rect 22190 8463 22246 8472
rect 22296 8430 22324 8842
rect 22284 8424 22336 8430
rect 22284 8366 22336 8372
rect 22388 8362 22416 9590
rect 22744 9580 22796 9586
rect 22744 9522 22796 9528
rect 22560 9376 22612 9382
rect 22560 9318 22612 9324
rect 22468 8832 22520 8838
rect 22468 8774 22520 8780
rect 22376 8356 22428 8362
rect 22376 8298 22428 8304
rect 22284 8288 22336 8294
rect 22284 8230 22336 8236
rect 22296 7886 22324 8230
rect 22284 7880 22336 7886
rect 22284 7822 22336 7828
rect 22112 6854 22232 6882
rect 22388 6866 22416 8298
rect 22480 7886 22508 8774
rect 22468 7880 22520 7886
rect 22468 7822 22520 7828
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 21836 6174 21956 6202
rect 21732 6112 21784 6118
rect 21732 6054 21784 6060
rect 21744 5914 21772 6054
rect 21732 5908 21784 5914
rect 21732 5850 21784 5856
rect 21836 5642 21864 6174
rect 21824 5636 21876 5642
rect 21824 5578 21876 5584
rect 21730 4720 21786 4729
rect 21730 4655 21732 4664
rect 21784 4655 21786 4664
rect 21732 4626 21784 4632
rect 21836 4026 21864 5578
rect 22008 5024 22060 5030
rect 22008 4966 22060 4972
rect 22020 4865 22048 4966
rect 22006 4856 22062 4865
rect 22006 4791 22008 4800
rect 22060 4791 22062 4800
rect 22008 4762 22060 4768
rect 22008 4616 22060 4622
rect 22008 4558 22060 4564
rect 22020 4282 22048 4558
rect 22008 4276 22060 4282
rect 22008 4218 22060 4224
rect 21744 4010 21864 4026
rect 21732 4004 21864 4010
rect 21784 3998 21864 4004
rect 21732 3946 21784 3952
rect 21836 2922 21864 3998
rect 22112 3942 22140 6734
rect 22204 6662 22232 6854
rect 22376 6860 22428 6866
rect 22376 6802 22428 6808
rect 22284 6792 22336 6798
rect 22284 6734 22336 6740
rect 22192 6656 22244 6662
rect 22192 6598 22244 6604
rect 22296 5574 22324 6734
rect 22480 6458 22508 7346
rect 22468 6452 22520 6458
rect 22468 6394 22520 6400
rect 22468 6248 22520 6254
rect 22468 6190 22520 6196
rect 22284 5568 22336 5574
rect 22284 5510 22336 5516
rect 22192 5364 22244 5370
rect 22192 5306 22244 5312
rect 22204 4690 22232 5306
rect 22480 4706 22508 6190
rect 22572 5710 22600 9318
rect 22652 8832 22704 8838
rect 22652 8774 22704 8780
rect 22664 8498 22692 8774
rect 22652 8492 22704 8498
rect 22652 8434 22704 8440
rect 22756 8090 22784 9522
rect 22848 9382 22876 9646
rect 22836 9376 22888 9382
rect 22836 9318 22888 9324
rect 22848 9042 22876 9318
rect 22836 9036 22888 9042
rect 22836 8978 22888 8984
rect 22744 8084 22796 8090
rect 22744 8026 22796 8032
rect 22836 6724 22888 6730
rect 22836 6666 22888 6672
rect 22848 6458 22876 6666
rect 22836 6452 22888 6458
rect 22836 6394 22888 6400
rect 22940 6390 22968 26318
rect 23020 24744 23072 24750
rect 23020 24686 23072 24692
rect 23032 21570 23060 24686
rect 23204 24268 23256 24274
rect 23204 24210 23256 24216
rect 23112 23520 23164 23526
rect 23112 23462 23164 23468
rect 23124 21690 23152 23462
rect 23112 21684 23164 21690
rect 23112 21626 23164 21632
rect 23032 21542 23152 21570
rect 23020 19712 23072 19718
rect 23020 19654 23072 19660
rect 23032 19446 23060 19654
rect 23020 19440 23072 19446
rect 23020 19382 23072 19388
rect 23124 18986 23152 21542
rect 23216 19922 23244 24210
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 23308 21026 23336 23802
rect 23388 23112 23440 23118
rect 23388 23054 23440 23060
rect 23400 21554 23428 23054
rect 23480 23044 23532 23050
rect 23480 22986 23532 22992
rect 23492 22778 23520 22986
rect 23480 22772 23532 22778
rect 23480 22714 23532 22720
rect 23492 22642 23520 22714
rect 23480 22636 23532 22642
rect 23480 22578 23532 22584
rect 23676 22094 23704 31232
rect 23756 29640 23808 29646
rect 23756 29582 23808 29588
rect 23768 29510 23796 29582
rect 23756 29504 23808 29510
rect 23756 29446 23808 29452
rect 23768 28937 23796 29446
rect 23848 29164 23900 29170
rect 23848 29106 23900 29112
rect 23754 28928 23810 28937
rect 23754 28863 23810 28872
rect 23860 28064 23888 29106
rect 23768 28036 23888 28064
rect 23768 26450 23796 28036
rect 23848 27940 23900 27946
rect 23848 27882 23900 27888
rect 23860 27606 23888 27882
rect 23848 27600 23900 27606
rect 23848 27542 23900 27548
rect 23860 27130 23888 27542
rect 23848 27124 23900 27130
rect 23848 27066 23900 27072
rect 23756 26444 23808 26450
rect 23756 26386 23808 26392
rect 23756 24064 23808 24070
rect 23756 24006 23808 24012
rect 23768 23186 23796 24006
rect 23756 23180 23808 23186
rect 23756 23122 23808 23128
rect 23952 22778 23980 34478
rect 24504 34105 24532 35430
rect 24490 34096 24546 34105
rect 24490 34031 24546 34040
rect 24768 33924 24820 33930
rect 24768 33866 24820 33872
rect 24032 33856 24084 33862
rect 24032 33798 24084 33804
rect 24044 32230 24072 33798
rect 24124 33516 24176 33522
rect 24124 33458 24176 33464
rect 24584 33516 24636 33522
rect 24584 33458 24636 33464
rect 24136 32434 24164 33458
rect 24596 32434 24624 33458
rect 24124 32428 24176 32434
rect 24124 32370 24176 32376
rect 24400 32428 24452 32434
rect 24400 32370 24452 32376
rect 24584 32428 24636 32434
rect 24584 32370 24636 32376
rect 24032 32224 24084 32230
rect 24032 32166 24084 32172
rect 24032 32020 24084 32026
rect 24032 31962 24084 31968
rect 24044 27674 24072 31962
rect 24124 31748 24176 31754
rect 24124 31690 24176 31696
rect 24136 30598 24164 31690
rect 24412 31686 24440 32370
rect 24400 31680 24452 31686
rect 24400 31622 24452 31628
rect 24216 31408 24268 31414
rect 24216 31350 24268 31356
rect 24228 30598 24256 31350
rect 24124 30592 24176 30598
rect 24124 30534 24176 30540
rect 24216 30592 24268 30598
rect 24216 30534 24268 30540
rect 24032 27668 24084 27674
rect 24032 27610 24084 27616
rect 24044 27402 24072 27610
rect 24032 27396 24084 27402
rect 24032 27338 24084 27344
rect 24032 26988 24084 26994
rect 24032 26930 24084 26936
rect 24044 26518 24072 26930
rect 24032 26512 24084 26518
rect 24032 26454 24084 26460
rect 24032 25220 24084 25226
rect 24032 25162 24084 25168
rect 24044 24954 24072 25162
rect 24032 24948 24084 24954
rect 24032 24890 24084 24896
rect 23940 22772 23992 22778
rect 23940 22714 23992 22720
rect 23848 22636 23900 22642
rect 23848 22578 23900 22584
rect 23756 22568 23808 22574
rect 23756 22510 23808 22516
rect 23584 22066 23704 22094
rect 23388 21548 23440 21554
rect 23388 21490 23440 21496
rect 23308 20998 23428 21026
rect 23296 20868 23348 20874
rect 23296 20810 23348 20816
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 23032 18958 23152 18986
rect 23032 14550 23060 18958
rect 23112 18896 23164 18902
rect 23112 18838 23164 18844
rect 23124 18358 23152 18838
rect 23308 18766 23336 20810
rect 23400 20058 23428 20998
rect 23584 20534 23612 22066
rect 23662 21992 23718 22001
rect 23662 21927 23718 21936
rect 23676 21622 23704 21927
rect 23664 21616 23716 21622
rect 23664 21558 23716 21564
rect 23664 21480 23716 21486
rect 23664 21422 23716 21428
rect 23676 21146 23704 21422
rect 23664 21140 23716 21146
rect 23664 21082 23716 21088
rect 23572 20528 23624 20534
rect 23572 20470 23624 20476
rect 23768 20262 23796 22510
rect 23860 21894 23888 22578
rect 23940 22092 23992 22098
rect 24136 22094 24164 30534
rect 24492 30320 24544 30326
rect 24492 30262 24544 30268
rect 24308 29708 24360 29714
rect 24308 29650 24360 29656
rect 24216 29640 24268 29646
rect 24216 29582 24268 29588
rect 24228 28422 24256 29582
rect 24320 29238 24348 29650
rect 24308 29232 24360 29238
rect 24308 29174 24360 29180
rect 24504 29170 24532 30262
rect 24596 29850 24624 32370
rect 24584 29844 24636 29850
rect 24584 29786 24636 29792
rect 24596 29306 24624 29786
rect 24780 29782 24808 33866
rect 24768 29776 24820 29782
rect 24768 29718 24820 29724
rect 24676 29640 24728 29646
rect 24676 29582 24728 29588
rect 24688 29510 24716 29582
rect 24676 29504 24728 29510
rect 24676 29446 24728 29452
rect 24584 29300 24636 29306
rect 24584 29242 24636 29248
rect 24492 29164 24544 29170
rect 24492 29106 24544 29112
rect 24216 28416 24268 28422
rect 24492 28416 24544 28422
rect 24216 28358 24268 28364
rect 24412 28376 24492 28404
rect 24216 28144 24268 28150
rect 24216 28086 24268 28092
rect 24228 27130 24256 28086
rect 24308 27872 24360 27878
rect 24308 27814 24360 27820
rect 24320 27713 24348 27814
rect 24306 27704 24362 27713
rect 24306 27639 24362 27648
rect 24412 27402 24440 28376
rect 24492 28358 24544 28364
rect 24400 27396 24452 27402
rect 24400 27338 24452 27344
rect 24216 27124 24268 27130
rect 24216 27066 24268 27072
rect 24216 26988 24268 26994
rect 24216 26930 24268 26936
rect 24228 25158 24256 26930
rect 24216 25152 24268 25158
rect 24216 25094 24268 25100
rect 24308 24336 24360 24342
rect 24308 24278 24360 24284
rect 24320 23798 24348 24278
rect 24308 23792 24360 23798
rect 24308 23734 24360 23740
rect 24412 23594 24440 27338
rect 24596 25770 24624 29242
rect 24676 29164 24728 29170
rect 24676 29106 24728 29112
rect 24584 25764 24636 25770
rect 24584 25706 24636 25712
rect 24688 25242 24716 29106
rect 24768 28416 24820 28422
rect 24768 28358 24820 28364
rect 24780 27946 24808 28358
rect 24768 27940 24820 27946
rect 24768 27882 24820 27888
rect 24872 26042 24900 39306
rect 25044 38752 25096 38758
rect 25044 38694 25096 38700
rect 25056 37262 25084 38694
rect 25148 38486 25176 39510
rect 25320 38752 25372 38758
rect 25320 38694 25372 38700
rect 25136 38480 25188 38486
rect 25332 38457 25360 38694
rect 25136 38422 25188 38428
rect 25318 38448 25374 38457
rect 25148 38010 25176 38422
rect 25318 38383 25374 38392
rect 25136 38004 25188 38010
rect 25136 37946 25188 37952
rect 25228 37868 25280 37874
rect 25148 37828 25228 37856
rect 25044 37256 25096 37262
rect 25044 37198 25096 37204
rect 25056 36786 25084 37198
rect 25044 36780 25096 36786
rect 25044 36722 25096 36728
rect 25044 35760 25096 35766
rect 25044 35702 25096 35708
rect 25056 33862 25084 35702
rect 25044 33856 25096 33862
rect 25044 33798 25096 33804
rect 25056 33522 25084 33798
rect 25044 33516 25096 33522
rect 25044 33458 25096 33464
rect 25056 32910 25084 33458
rect 25044 32904 25096 32910
rect 25044 32846 25096 32852
rect 25056 31346 25084 32846
rect 25044 31340 25096 31346
rect 25044 31282 25096 31288
rect 25044 30728 25096 30734
rect 25044 30670 25096 30676
rect 24952 30388 25004 30394
rect 24952 30330 25004 30336
rect 24964 29617 24992 30330
rect 25056 29730 25084 30670
rect 25148 30394 25176 37828
rect 25228 37810 25280 37816
rect 25320 37188 25372 37194
rect 25320 37130 25372 37136
rect 25332 34950 25360 37130
rect 25516 36106 25544 40054
rect 25964 39364 26016 39370
rect 25964 39306 26016 39312
rect 25504 36100 25556 36106
rect 25504 36042 25556 36048
rect 25976 36038 26004 39306
rect 26240 39296 26292 39302
rect 26240 39238 26292 39244
rect 26252 38554 26280 39238
rect 26424 38956 26476 38962
rect 26424 38898 26476 38904
rect 26240 38548 26292 38554
rect 26240 38490 26292 38496
rect 26436 38486 26464 38898
rect 26424 38480 26476 38486
rect 26424 38422 26476 38428
rect 26056 38344 26108 38350
rect 26056 38286 26108 38292
rect 26332 38344 26384 38350
rect 26332 38286 26384 38292
rect 26068 37806 26096 38286
rect 26344 37874 26372 38286
rect 26332 37868 26384 37874
rect 26332 37810 26384 37816
rect 26056 37800 26108 37806
rect 26056 37742 26108 37748
rect 25688 36032 25740 36038
rect 25688 35974 25740 35980
rect 25872 36032 25924 36038
rect 25872 35974 25924 35980
rect 25964 36032 26016 36038
rect 25964 35974 26016 35980
rect 25504 35556 25556 35562
rect 25504 35498 25556 35504
rect 25516 35222 25544 35498
rect 25504 35216 25556 35222
rect 25504 35158 25556 35164
rect 25700 35018 25728 35974
rect 25780 35760 25832 35766
rect 25780 35702 25832 35708
rect 25688 35012 25740 35018
rect 25688 34954 25740 34960
rect 25320 34944 25372 34950
rect 25320 34886 25372 34892
rect 25320 32836 25372 32842
rect 25320 32778 25372 32784
rect 25332 32570 25360 32778
rect 25320 32564 25372 32570
rect 25320 32506 25372 32512
rect 25596 32428 25648 32434
rect 25596 32370 25648 32376
rect 25320 32360 25372 32366
rect 25320 32302 25372 32308
rect 25228 31340 25280 31346
rect 25228 31282 25280 31288
rect 25240 30938 25268 31282
rect 25228 30932 25280 30938
rect 25228 30874 25280 30880
rect 25136 30388 25188 30394
rect 25136 30330 25188 30336
rect 25056 29702 25176 29730
rect 25044 29640 25096 29646
rect 24950 29608 25006 29617
rect 25044 29582 25096 29588
rect 24950 29543 25006 29552
rect 24860 26036 24912 26042
rect 24860 25978 24912 25984
rect 24688 25226 24900 25242
rect 24688 25220 24912 25226
rect 24688 25214 24860 25220
rect 24860 25162 24912 25168
rect 24768 25152 24820 25158
rect 24768 25094 24820 25100
rect 24492 24812 24544 24818
rect 24492 24754 24544 24760
rect 24676 24812 24728 24818
rect 24676 24754 24728 24760
rect 24504 24410 24532 24754
rect 24492 24404 24544 24410
rect 24492 24346 24544 24352
rect 24688 23905 24716 24754
rect 24674 23896 24730 23905
rect 24674 23831 24730 23840
rect 24400 23588 24452 23594
rect 24400 23530 24452 23536
rect 24136 22066 24256 22094
rect 23940 22034 23992 22040
rect 23848 21888 23900 21894
rect 23848 21830 23900 21836
rect 23480 20256 23532 20262
rect 23480 20198 23532 20204
rect 23756 20256 23808 20262
rect 23756 20198 23808 20204
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 23492 19854 23520 20198
rect 23572 19916 23624 19922
rect 23572 19858 23624 19864
rect 23480 19848 23532 19854
rect 23480 19790 23532 19796
rect 23584 18834 23612 19858
rect 23756 19780 23808 19786
rect 23756 19722 23808 19728
rect 23768 19378 23796 19722
rect 23756 19372 23808 19378
rect 23756 19314 23808 19320
rect 23572 18828 23624 18834
rect 23572 18770 23624 18776
rect 23296 18760 23348 18766
rect 23296 18702 23348 18708
rect 23204 18692 23256 18698
rect 23204 18634 23256 18640
rect 23112 18352 23164 18358
rect 23112 18294 23164 18300
rect 23216 18068 23244 18634
rect 23388 18624 23440 18630
rect 23388 18566 23440 18572
rect 23400 18290 23428 18566
rect 23388 18284 23440 18290
rect 23388 18226 23440 18232
rect 23296 18080 23348 18086
rect 23216 18040 23296 18068
rect 23216 17678 23244 18040
rect 23296 18022 23348 18028
rect 23296 17876 23348 17882
rect 23296 17818 23348 17824
rect 23204 17672 23256 17678
rect 23204 17614 23256 17620
rect 23308 17202 23336 17818
rect 23296 17196 23348 17202
rect 23296 17138 23348 17144
rect 23308 17105 23336 17138
rect 23294 17096 23350 17105
rect 23294 17031 23350 17040
rect 23400 16522 23428 18226
rect 23480 16584 23532 16590
rect 23480 16526 23532 16532
rect 23296 16516 23348 16522
rect 23296 16458 23348 16464
rect 23388 16516 23440 16522
rect 23388 16458 23440 16464
rect 23112 16448 23164 16454
rect 23112 16390 23164 16396
rect 23124 16182 23152 16390
rect 23112 16176 23164 16182
rect 23112 16118 23164 16124
rect 23308 15706 23336 16458
rect 23492 16250 23520 16526
rect 23480 16244 23532 16250
rect 23480 16186 23532 16192
rect 23848 16176 23900 16182
rect 23848 16118 23900 16124
rect 23480 15904 23532 15910
rect 23480 15846 23532 15852
rect 23296 15700 23348 15706
rect 23296 15642 23348 15648
rect 23492 15502 23520 15846
rect 23480 15496 23532 15502
rect 23480 15438 23532 15444
rect 23860 15026 23888 16118
rect 23848 15020 23900 15026
rect 23848 14962 23900 14968
rect 23020 14544 23072 14550
rect 23020 14486 23072 14492
rect 23952 14346 23980 22034
rect 24032 21548 24084 21554
rect 24032 21490 24084 21496
rect 24044 19514 24072 21490
rect 24124 20392 24176 20398
rect 24124 20334 24176 20340
rect 24032 19508 24084 19514
rect 24032 19450 24084 19456
rect 24136 18290 24164 20334
rect 24124 18284 24176 18290
rect 24124 18226 24176 18232
rect 23940 14340 23992 14346
rect 23940 14282 23992 14288
rect 23112 14272 23164 14278
rect 23112 14214 23164 14220
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 23032 11354 23060 12242
rect 23020 11348 23072 11354
rect 23020 11290 23072 11296
rect 23124 11234 23152 14214
rect 23664 13932 23716 13938
rect 23664 13874 23716 13880
rect 23676 13530 23704 13874
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 23756 13252 23808 13258
rect 23756 13194 23808 13200
rect 23768 12850 23796 13194
rect 23756 12844 23808 12850
rect 23756 12786 23808 12792
rect 23480 12640 23532 12646
rect 23480 12582 23532 12588
rect 23664 12640 23716 12646
rect 23664 12582 23716 12588
rect 23492 12442 23520 12582
rect 23480 12436 23532 12442
rect 23480 12378 23532 12384
rect 23480 12232 23532 12238
rect 23480 12174 23532 12180
rect 23492 11286 23520 12174
rect 23032 11206 23152 11234
rect 23480 11280 23532 11286
rect 23480 11222 23532 11228
rect 23032 11150 23060 11206
rect 23020 11144 23072 11150
rect 23020 11086 23072 11092
rect 23032 10062 23060 11086
rect 23020 10056 23072 10062
rect 23020 9998 23072 10004
rect 23204 9648 23256 9654
rect 23204 9590 23256 9596
rect 23112 9512 23164 9518
rect 23112 9454 23164 9460
rect 23020 8968 23072 8974
rect 23020 8910 23072 8916
rect 23032 7410 23060 8910
rect 23124 8294 23152 9454
rect 23216 8974 23244 9590
rect 23204 8968 23256 8974
rect 23204 8910 23256 8916
rect 23112 8288 23164 8294
rect 23112 8230 23164 8236
rect 23216 7886 23244 8910
rect 23296 8560 23348 8566
rect 23296 8502 23348 8508
rect 23480 8560 23532 8566
rect 23480 8502 23532 8508
rect 23308 7954 23336 8502
rect 23296 7948 23348 7954
rect 23296 7890 23348 7896
rect 23204 7880 23256 7886
rect 23204 7822 23256 7828
rect 23020 7404 23072 7410
rect 23020 7346 23072 7352
rect 23020 7200 23072 7206
rect 23020 7142 23072 7148
rect 22928 6384 22980 6390
rect 22928 6326 22980 6332
rect 23032 6322 23060 7142
rect 23020 6316 23072 6322
rect 23020 6258 23072 6264
rect 22744 6248 22796 6254
rect 22744 6190 22796 6196
rect 22560 5704 22612 5710
rect 22560 5646 22612 5652
rect 22572 5302 22600 5646
rect 22560 5296 22612 5302
rect 22560 5238 22612 5244
rect 22192 4684 22244 4690
rect 22480 4678 22600 4706
rect 22192 4626 22244 4632
rect 22468 4616 22520 4622
rect 22468 4558 22520 4564
rect 22192 4480 22244 4486
rect 22192 4422 22244 4428
rect 22284 4480 22336 4486
rect 22284 4422 22336 4428
rect 22204 4214 22232 4422
rect 22192 4208 22244 4214
rect 22192 4150 22244 4156
rect 22100 3936 22152 3942
rect 22100 3878 22152 3884
rect 22112 3602 22140 3878
rect 22100 3596 22152 3602
rect 22100 3538 22152 3544
rect 22296 2938 22324 4422
rect 22480 3194 22508 4558
rect 22572 3942 22600 4678
rect 22560 3936 22612 3942
rect 22560 3878 22612 3884
rect 22468 3188 22520 3194
rect 22468 3130 22520 3136
rect 22376 3052 22428 3058
rect 22376 2994 22428 3000
rect 21824 2916 21876 2922
rect 21824 2858 21876 2864
rect 22020 2910 22324 2938
rect 22020 800 22048 2910
rect 22388 800 22416 2994
rect 22756 800 22784 6190
rect 23216 5234 23244 7822
rect 23492 7818 23520 8502
rect 23296 7812 23348 7818
rect 23296 7754 23348 7760
rect 23480 7812 23532 7818
rect 23480 7754 23532 7760
rect 23308 6730 23336 7754
rect 23492 7478 23520 7754
rect 23572 7744 23624 7750
rect 23572 7686 23624 7692
rect 23480 7472 23532 7478
rect 23480 7414 23532 7420
rect 23296 6724 23348 6730
rect 23296 6666 23348 6672
rect 23584 5778 23612 7686
rect 23572 5772 23624 5778
rect 23572 5714 23624 5720
rect 23204 5228 23256 5234
rect 23204 5170 23256 5176
rect 23216 5030 23244 5170
rect 23204 5024 23256 5030
rect 23204 4966 23256 4972
rect 23676 4622 23704 12582
rect 23952 7410 23980 14282
rect 24124 12232 24176 12238
rect 24124 12174 24176 12180
rect 24032 12096 24084 12102
rect 24032 12038 24084 12044
rect 24044 11830 24072 12038
rect 24136 11830 24164 12174
rect 24032 11824 24084 11830
rect 24032 11766 24084 11772
rect 24124 11824 24176 11830
rect 24124 11766 24176 11772
rect 24136 11218 24164 11766
rect 24124 11212 24176 11218
rect 24124 11154 24176 11160
rect 24228 8498 24256 22066
rect 24780 22030 24808 25094
rect 24872 24886 24900 25162
rect 24860 24880 24912 24886
rect 24860 24822 24912 24828
rect 24872 24206 24900 24822
rect 24860 24200 24912 24206
rect 24860 24142 24912 24148
rect 24964 22030 24992 29543
rect 25056 28082 25084 29582
rect 25148 29073 25176 29702
rect 25134 29064 25190 29073
rect 25134 28999 25190 29008
rect 25044 28076 25096 28082
rect 25044 28018 25096 28024
rect 25148 24682 25176 28999
rect 25332 28234 25360 32302
rect 25608 32026 25636 32370
rect 25596 32020 25648 32026
rect 25596 31962 25648 31968
rect 25700 31754 25728 34954
rect 25792 34746 25820 35702
rect 25884 35494 25912 35974
rect 25872 35488 25924 35494
rect 25872 35430 25924 35436
rect 25964 35080 26016 35086
rect 25964 35022 26016 35028
rect 25780 34740 25832 34746
rect 25780 34682 25832 34688
rect 25976 34542 26004 35022
rect 25964 34536 26016 34542
rect 25964 34478 26016 34484
rect 25778 32872 25834 32881
rect 25778 32807 25834 32816
rect 25792 32570 25820 32807
rect 25780 32564 25832 32570
rect 25780 32506 25832 32512
rect 25792 32434 25820 32506
rect 25780 32428 25832 32434
rect 25780 32370 25832 32376
rect 25872 32292 25924 32298
rect 25872 32234 25924 32240
rect 25884 31890 25912 32234
rect 25872 31884 25924 31890
rect 25872 31826 25924 31832
rect 25608 31726 25728 31754
rect 26068 31754 26096 37742
rect 27264 37262 27292 41482
rect 27724 38010 27752 42706
rect 27988 41540 28040 41546
rect 27988 41482 28040 41488
rect 27712 38004 27764 38010
rect 27712 37946 27764 37952
rect 27896 37936 27948 37942
rect 27896 37878 27948 37884
rect 27252 37256 27304 37262
rect 26422 37224 26478 37233
rect 27252 37198 27304 37204
rect 26422 37159 26478 37168
rect 26436 36922 26464 37159
rect 26792 37120 26844 37126
rect 26792 37062 26844 37068
rect 26424 36916 26476 36922
rect 26424 36858 26476 36864
rect 26804 36854 26832 37062
rect 26792 36848 26844 36854
rect 26792 36790 26844 36796
rect 26332 36780 26384 36786
rect 26332 36722 26384 36728
rect 26344 36310 26372 36722
rect 26332 36304 26384 36310
rect 26332 36246 26384 36252
rect 26516 36168 26568 36174
rect 26516 36110 26568 36116
rect 26528 35834 26556 36110
rect 26516 35828 26568 35834
rect 26516 35770 26568 35776
rect 26332 35080 26384 35086
rect 26332 35022 26384 35028
rect 26344 34610 26372 35022
rect 26332 34604 26384 34610
rect 26332 34546 26384 34552
rect 26148 34536 26200 34542
rect 26148 34478 26200 34484
rect 26160 32774 26188 34478
rect 26148 32768 26200 32774
rect 26148 32710 26200 32716
rect 26160 32366 26188 32710
rect 26148 32360 26200 32366
rect 26148 32302 26200 32308
rect 26068 31726 26188 31754
rect 25412 31680 25464 31686
rect 25412 31622 25464 31628
rect 25424 30870 25452 31622
rect 25412 30864 25464 30870
rect 25412 30806 25464 30812
rect 25608 28642 25636 31726
rect 26160 31142 26188 31726
rect 26148 31136 26200 31142
rect 26148 31078 26200 31084
rect 26160 30802 26188 31078
rect 26148 30796 26200 30802
rect 26148 30738 26200 30744
rect 25872 30728 25924 30734
rect 25872 30670 25924 30676
rect 25884 30122 25912 30670
rect 25872 30116 25924 30122
rect 25872 30058 25924 30064
rect 25780 30048 25832 30054
rect 25780 29990 25832 29996
rect 25688 29572 25740 29578
rect 25688 29514 25740 29520
rect 25700 29306 25728 29514
rect 25688 29300 25740 29306
rect 25688 29242 25740 29248
rect 25792 29170 25820 29990
rect 25780 29164 25832 29170
rect 25780 29106 25832 29112
rect 25872 29164 25924 29170
rect 26056 29164 26108 29170
rect 25872 29106 25924 29112
rect 25976 29124 26056 29152
rect 25792 29034 25820 29106
rect 25780 29028 25832 29034
rect 25780 28970 25832 28976
rect 25884 28762 25912 29106
rect 25976 29034 26004 29124
rect 26056 29106 26108 29112
rect 25964 29028 26016 29034
rect 25964 28970 26016 28976
rect 25872 28756 25924 28762
rect 25872 28698 25924 28704
rect 25240 28206 25360 28234
rect 25424 28614 25636 28642
rect 25136 24676 25188 24682
rect 25136 24618 25188 24624
rect 25044 24200 25096 24206
rect 25044 24142 25096 24148
rect 25056 23730 25084 24142
rect 25136 23860 25188 23866
rect 25136 23802 25188 23808
rect 25044 23724 25096 23730
rect 25044 23666 25096 23672
rect 25056 23118 25084 23666
rect 25044 23112 25096 23118
rect 25044 23054 25096 23060
rect 25148 22642 25176 23802
rect 25044 22636 25096 22642
rect 25044 22578 25096 22584
rect 25136 22636 25188 22642
rect 25136 22578 25188 22584
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 24952 22024 25004 22030
rect 24952 21966 25004 21972
rect 24584 21888 24636 21894
rect 24584 21830 24636 21836
rect 24596 21418 24624 21830
rect 25056 21690 25084 22578
rect 25136 22024 25188 22030
rect 25136 21966 25188 21972
rect 25148 21865 25176 21966
rect 25134 21856 25190 21865
rect 25134 21791 25190 21800
rect 25044 21684 25096 21690
rect 25044 21626 25096 21632
rect 24584 21412 24636 21418
rect 24584 21354 24636 21360
rect 24400 21344 24452 21350
rect 24400 21286 24452 21292
rect 24412 20942 24440 21286
rect 24596 20942 24624 21354
rect 24676 21072 24728 21078
rect 24676 21014 24728 21020
rect 24400 20936 24452 20942
rect 24400 20878 24452 20884
rect 24584 20936 24636 20942
rect 24584 20878 24636 20884
rect 24688 20874 24716 21014
rect 24308 20868 24360 20874
rect 24308 20810 24360 20816
rect 24676 20868 24728 20874
rect 24676 20810 24728 20816
rect 24320 20398 24348 20810
rect 24584 20800 24636 20806
rect 24584 20742 24636 20748
rect 24492 20460 24544 20466
rect 24492 20402 24544 20408
rect 24308 20392 24360 20398
rect 24308 20334 24360 20340
rect 24320 19174 24348 20334
rect 24504 19854 24532 20402
rect 24492 19848 24544 19854
rect 24492 19790 24544 19796
rect 24400 19372 24452 19378
rect 24400 19314 24452 19320
rect 24308 19168 24360 19174
rect 24308 19110 24360 19116
rect 24320 18358 24348 19110
rect 24412 18970 24440 19314
rect 24400 18964 24452 18970
rect 24400 18906 24452 18912
rect 24492 18692 24544 18698
rect 24492 18634 24544 18640
rect 24308 18352 24360 18358
rect 24308 18294 24360 18300
rect 24504 18154 24532 18634
rect 24492 18148 24544 18154
rect 24492 18090 24544 18096
rect 24596 16590 24624 20742
rect 24860 20392 24912 20398
rect 24860 20334 24912 20340
rect 24676 20256 24728 20262
rect 24676 20198 24728 20204
rect 24688 19922 24716 20198
rect 24676 19916 24728 19922
rect 24676 19858 24728 19864
rect 24872 19854 24900 20334
rect 24860 19848 24912 19854
rect 24860 19790 24912 19796
rect 24952 19712 25004 19718
rect 24766 19680 24822 19689
rect 24952 19654 25004 19660
rect 24766 19615 24822 19624
rect 24780 19514 24808 19615
rect 24768 19508 24820 19514
rect 24768 19450 24820 19456
rect 24676 18148 24728 18154
rect 24676 18090 24728 18096
rect 24688 17785 24716 18090
rect 24674 17776 24730 17785
rect 24674 17711 24730 17720
rect 24676 17196 24728 17202
rect 24676 17138 24728 17144
rect 24584 16584 24636 16590
rect 24584 16526 24636 16532
rect 24400 16448 24452 16454
rect 24400 16390 24452 16396
rect 24412 16182 24440 16390
rect 24688 16250 24716 17138
rect 24676 16244 24728 16250
rect 24676 16186 24728 16192
rect 24400 16176 24452 16182
rect 24400 16118 24452 16124
rect 24492 15972 24544 15978
rect 24492 15914 24544 15920
rect 24308 14816 24360 14822
rect 24308 14758 24360 14764
rect 24216 8492 24268 8498
rect 24216 8434 24268 8440
rect 23940 7404 23992 7410
rect 23940 7346 23992 7352
rect 24124 6860 24176 6866
rect 24124 6802 24176 6808
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 23664 4616 23716 4622
rect 23664 4558 23716 4564
rect 23480 4480 23532 4486
rect 23480 4422 23532 4428
rect 23492 3618 23520 4422
rect 23124 3590 23520 3618
rect 23572 3596 23624 3602
rect 23124 800 23152 3590
rect 23572 3538 23624 3544
rect 23296 3528 23348 3534
rect 23296 3470 23348 3476
rect 23308 2650 23336 3470
rect 23584 3058 23612 3538
rect 23572 3052 23624 3058
rect 23572 2994 23624 3000
rect 23480 2848 23532 2854
rect 23480 2790 23532 2796
rect 23296 2644 23348 2650
rect 23296 2586 23348 2592
rect 23492 2446 23520 2790
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 23492 870 23612 898
rect 23492 800 23520 870
rect 19904 734 20116 762
rect 20166 0 20222 800
rect 20534 0 20590 800
rect 20902 0 20958 800
rect 21270 0 21326 800
rect 21638 0 21694 800
rect 22006 0 22062 800
rect 22374 0 22430 800
rect 22742 0 22798 800
rect 23110 0 23166 800
rect 23478 0 23534 800
rect 23584 762 23612 870
rect 23768 762 23796 6258
rect 23848 6112 23900 6118
rect 23848 6054 23900 6060
rect 23860 3126 23888 6054
rect 23940 5636 23992 5642
rect 23940 5578 23992 5584
rect 23952 4729 23980 5578
rect 23938 4720 23994 4729
rect 23938 4655 23940 4664
rect 23992 4655 23994 4664
rect 23940 4626 23992 4632
rect 23952 4595 23980 4626
rect 23848 3120 23900 3126
rect 23848 3062 23900 3068
rect 24136 2774 24164 6802
rect 23860 2746 24164 2774
rect 23860 800 23888 2746
rect 24320 2582 24348 14758
rect 24400 13728 24452 13734
rect 24400 13670 24452 13676
rect 24412 13326 24440 13670
rect 24504 13530 24532 15914
rect 24688 15502 24716 16186
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24780 14346 24808 19450
rect 24860 19440 24912 19446
rect 24860 19382 24912 19388
rect 24872 17746 24900 19382
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 24860 16040 24912 16046
rect 24860 15982 24912 15988
rect 24872 14618 24900 15982
rect 24860 14612 24912 14618
rect 24860 14554 24912 14560
rect 24768 14340 24820 14346
rect 24768 14282 24820 14288
rect 24780 14074 24808 14282
rect 24768 14068 24820 14074
rect 24768 14010 24820 14016
rect 24872 14006 24900 14554
rect 24860 14000 24912 14006
rect 24860 13942 24912 13948
rect 24492 13524 24544 13530
rect 24492 13466 24544 13472
rect 24964 13394 24992 19654
rect 25056 19446 25084 21626
rect 25136 21140 25188 21146
rect 25136 21082 25188 21088
rect 25148 21010 25176 21082
rect 25136 21004 25188 21010
rect 25136 20946 25188 20952
rect 25240 20466 25268 28206
rect 25320 28076 25372 28082
rect 25320 28018 25372 28024
rect 25332 27130 25360 28018
rect 25320 27124 25372 27130
rect 25320 27066 25372 27072
rect 25320 24132 25372 24138
rect 25320 24074 25372 24080
rect 25332 23730 25360 24074
rect 25320 23724 25372 23730
rect 25320 23666 25372 23672
rect 25320 21888 25372 21894
rect 25320 21830 25372 21836
rect 25332 21146 25360 21830
rect 25320 21140 25372 21146
rect 25320 21082 25372 21088
rect 25424 20602 25452 28614
rect 25596 28484 25648 28490
rect 25596 28426 25648 28432
rect 25608 26994 25636 28426
rect 26160 27470 26188 30738
rect 26344 28218 26372 34546
rect 26516 33924 26568 33930
rect 26516 33866 26568 33872
rect 26528 33658 26556 33866
rect 27264 33658 27292 37198
rect 27620 37188 27672 37194
rect 27620 37130 27672 37136
rect 27632 36922 27660 37130
rect 27620 36916 27672 36922
rect 27620 36858 27672 36864
rect 27908 36106 27936 37878
rect 27896 36100 27948 36106
rect 27896 36042 27948 36048
rect 27908 35766 27936 36042
rect 27896 35760 27948 35766
rect 27896 35702 27948 35708
rect 27804 35080 27856 35086
rect 27804 35022 27856 35028
rect 27816 34474 27844 35022
rect 28000 34746 28028 41482
rect 28184 37738 28212 47058
rect 29656 46578 29684 49286
rect 30378 49200 30434 50000
rect 31206 49314 31262 50000
rect 32034 49314 32090 50000
rect 31206 49286 31524 49314
rect 31206 49200 31262 49286
rect 29828 47048 29880 47054
rect 29828 46990 29880 46996
rect 29644 46572 29696 46578
rect 29644 46514 29696 46520
rect 28356 38004 28408 38010
rect 28356 37946 28408 37952
rect 28368 37806 28396 37946
rect 28356 37800 28408 37806
rect 28356 37742 28408 37748
rect 28172 37732 28224 37738
rect 28172 37674 28224 37680
rect 28264 35828 28316 35834
rect 28264 35770 28316 35776
rect 28172 35556 28224 35562
rect 28172 35498 28224 35504
rect 28184 35290 28212 35498
rect 28172 35284 28224 35290
rect 28172 35226 28224 35232
rect 28080 34944 28132 34950
rect 28080 34886 28132 34892
rect 27988 34740 28040 34746
rect 27988 34682 28040 34688
rect 27804 34468 27856 34474
rect 27804 34410 27856 34416
rect 28092 33998 28120 34886
rect 28276 34542 28304 35770
rect 28368 35578 28396 37742
rect 28540 37732 28592 37738
rect 28540 37674 28592 37680
rect 28552 36718 28580 37674
rect 29552 37664 29604 37670
rect 29552 37606 29604 37612
rect 28908 37324 28960 37330
rect 28908 37266 28960 37272
rect 28632 36848 28684 36854
rect 28632 36790 28684 36796
rect 28540 36712 28592 36718
rect 28540 36654 28592 36660
rect 28552 36242 28580 36654
rect 28540 36236 28592 36242
rect 28540 36178 28592 36184
rect 28448 36168 28500 36174
rect 28448 36110 28500 36116
rect 28460 35698 28488 36110
rect 28540 36032 28592 36038
rect 28540 35974 28592 35980
rect 28448 35692 28500 35698
rect 28448 35634 28500 35640
rect 28368 35550 28488 35578
rect 28552 35562 28580 35974
rect 28644 35834 28672 36790
rect 28816 36168 28868 36174
rect 28816 36110 28868 36116
rect 28632 35828 28684 35834
rect 28632 35770 28684 35776
rect 28828 35698 28856 36110
rect 28724 35692 28776 35698
rect 28724 35634 28776 35640
rect 28816 35692 28868 35698
rect 28816 35634 28868 35640
rect 28264 34536 28316 34542
rect 28264 34478 28316 34484
rect 28080 33992 28132 33998
rect 28080 33934 28132 33940
rect 27528 33856 27580 33862
rect 27528 33798 27580 33804
rect 27896 33856 27948 33862
rect 27896 33798 27948 33804
rect 26516 33652 26568 33658
rect 26516 33594 26568 33600
rect 27252 33652 27304 33658
rect 27252 33594 27304 33600
rect 27540 33522 27568 33798
rect 27908 33590 27936 33798
rect 27896 33584 27948 33590
rect 27896 33526 27948 33532
rect 27528 33516 27580 33522
rect 27528 33458 27580 33464
rect 27804 33516 27856 33522
rect 27804 33458 27856 33464
rect 27620 32904 27672 32910
rect 27620 32846 27672 32852
rect 27436 32428 27488 32434
rect 27436 32370 27488 32376
rect 27448 32026 27476 32370
rect 27436 32020 27488 32026
rect 27436 31962 27488 31968
rect 27528 31680 27580 31686
rect 27528 31622 27580 31628
rect 27540 31482 27568 31622
rect 27528 31476 27580 31482
rect 27528 31418 27580 31424
rect 27632 29730 27660 32846
rect 27712 32564 27764 32570
rect 27712 32506 27764 32512
rect 27724 32434 27752 32506
rect 27712 32428 27764 32434
rect 27712 32370 27764 32376
rect 27816 32230 27844 33458
rect 28172 32836 28224 32842
rect 28172 32778 28224 32784
rect 28184 32570 28212 32778
rect 28172 32564 28224 32570
rect 28172 32506 28224 32512
rect 28276 32450 28304 34478
rect 28184 32422 28304 32450
rect 28356 32428 28408 32434
rect 27804 32224 27856 32230
rect 27804 32166 27856 32172
rect 27804 31884 27856 31890
rect 27804 31826 27856 31832
rect 27712 30592 27764 30598
rect 27712 30534 27764 30540
rect 27540 29714 27660 29730
rect 27528 29708 27660 29714
rect 27580 29702 27660 29708
rect 27528 29650 27580 29656
rect 26976 29504 27028 29510
rect 26976 29446 27028 29452
rect 26988 28490 27016 29446
rect 27528 28960 27580 28966
rect 27528 28902 27580 28908
rect 27540 28694 27568 28902
rect 27528 28688 27580 28694
rect 27528 28630 27580 28636
rect 26976 28484 27028 28490
rect 26976 28426 27028 28432
rect 26792 28416 26844 28422
rect 26792 28358 26844 28364
rect 26332 28212 26384 28218
rect 26332 28154 26384 28160
rect 25872 27464 25924 27470
rect 25872 27406 25924 27412
rect 26148 27464 26200 27470
rect 26148 27406 26200 27412
rect 26240 27464 26292 27470
rect 26344 27452 26372 28154
rect 26804 27674 26832 28358
rect 26988 28082 27016 28426
rect 26976 28076 27028 28082
rect 26976 28018 27028 28024
rect 26988 27690 27016 28018
rect 27632 27878 27660 29702
rect 27724 29306 27752 30534
rect 27816 30394 27844 31826
rect 27988 31816 28040 31822
rect 27988 31758 28040 31764
rect 28000 31346 28028 31758
rect 27988 31340 28040 31346
rect 27988 31282 28040 31288
rect 27988 31204 28040 31210
rect 27988 31146 28040 31152
rect 27804 30388 27856 30394
rect 27804 30330 27856 30336
rect 27804 29572 27856 29578
rect 27804 29514 27856 29520
rect 27712 29300 27764 29306
rect 27712 29242 27764 29248
rect 27816 28762 27844 29514
rect 27896 28960 27948 28966
rect 27896 28902 27948 28908
rect 27804 28756 27856 28762
rect 27804 28698 27856 28704
rect 27908 28558 27936 28902
rect 27896 28552 27948 28558
rect 27896 28494 27948 28500
rect 28000 28422 28028 31146
rect 28080 30592 28132 30598
rect 28080 30534 28132 30540
rect 28092 30258 28120 30534
rect 28080 30252 28132 30258
rect 28080 30194 28132 30200
rect 28080 30116 28132 30122
rect 28080 30058 28132 30064
rect 28092 29073 28120 30058
rect 28078 29064 28134 29073
rect 28078 28999 28134 29008
rect 28092 28558 28120 28999
rect 28080 28552 28132 28558
rect 28080 28494 28132 28500
rect 27988 28416 28040 28422
rect 27988 28358 28040 28364
rect 27620 27872 27672 27878
rect 27620 27814 27672 27820
rect 26792 27668 26844 27674
rect 26988 27662 27200 27690
rect 26792 27610 26844 27616
rect 26424 27464 26476 27470
rect 26344 27424 26424 27452
rect 26240 27406 26292 27412
rect 26424 27406 26476 27412
rect 25884 27130 25912 27406
rect 25872 27124 25924 27130
rect 25872 27066 25924 27072
rect 25596 26988 25648 26994
rect 25596 26930 25648 26936
rect 25504 26920 25556 26926
rect 25504 26862 25556 26868
rect 25516 26314 25544 26862
rect 25504 26308 25556 26314
rect 25504 26250 25556 26256
rect 25504 23724 25556 23730
rect 25504 23666 25556 23672
rect 25516 23322 25544 23666
rect 25504 23316 25556 23322
rect 25504 23258 25556 23264
rect 25608 22094 25636 26930
rect 26252 26790 26280 27406
rect 26240 26784 26292 26790
rect 26240 26726 26292 26732
rect 26252 26586 26280 26726
rect 26240 26580 26292 26586
rect 26240 26522 26292 26528
rect 26240 26036 26292 26042
rect 26240 25978 26292 25984
rect 25688 25900 25740 25906
rect 26056 25900 26108 25906
rect 25740 25860 25820 25888
rect 25688 25842 25740 25848
rect 25792 25158 25820 25860
rect 26056 25842 26108 25848
rect 25964 25832 26016 25838
rect 25964 25774 26016 25780
rect 25976 25362 26004 25774
rect 25964 25356 26016 25362
rect 25964 25298 26016 25304
rect 25780 25152 25832 25158
rect 25780 25094 25832 25100
rect 25792 24954 25820 25094
rect 25780 24948 25832 24954
rect 25780 24890 25832 24896
rect 25686 24168 25742 24177
rect 25686 24103 25742 24112
rect 25700 24070 25728 24103
rect 25688 24064 25740 24070
rect 25688 24006 25740 24012
rect 25700 23730 25728 24006
rect 25792 23866 25820 24890
rect 25964 24812 26016 24818
rect 25964 24754 26016 24760
rect 25976 24614 26004 24754
rect 25964 24608 26016 24614
rect 25964 24550 26016 24556
rect 25976 24342 26004 24550
rect 25964 24336 26016 24342
rect 25964 24278 26016 24284
rect 26068 24018 26096 25842
rect 26148 24132 26200 24138
rect 26148 24074 26200 24080
rect 25884 23990 26096 24018
rect 25780 23860 25832 23866
rect 25780 23802 25832 23808
rect 25884 23746 25912 23990
rect 26056 23860 26108 23866
rect 26056 23802 26108 23808
rect 25688 23724 25740 23730
rect 25688 23666 25740 23672
rect 25792 23718 25912 23746
rect 25792 23168 25820 23718
rect 25872 23656 25924 23662
rect 25872 23598 25924 23604
rect 25516 22066 25636 22094
rect 25700 23140 25820 23168
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25410 20496 25466 20505
rect 25136 20460 25188 20466
rect 25136 20402 25188 20408
rect 25228 20460 25280 20466
rect 25410 20431 25412 20440
rect 25228 20402 25280 20408
rect 25464 20431 25466 20440
rect 25412 20402 25464 20408
rect 25148 19990 25176 20402
rect 25228 20052 25280 20058
rect 25228 19994 25280 20000
rect 25136 19984 25188 19990
rect 25136 19926 25188 19932
rect 25148 19854 25176 19926
rect 25136 19848 25188 19854
rect 25136 19790 25188 19796
rect 25044 19440 25096 19446
rect 25044 19382 25096 19388
rect 25044 18352 25096 18358
rect 25044 18294 25096 18300
rect 25056 17066 25084 18294
rect 25148 18086 25176 19790
rect 25240 18766 25268 19994
rect 25424 19786 25452 20402
rect 25412 19780 25464 19786
rect 25412 19722 25464 19728
rect 25228 18760 25280 18766
rect 25228 18702 25280 18708
rect 25228 18624 25280 18630
rect 25228 18566 25280 18572
rect 25136 18080 25188 18086
rect 25136 18022 25188 18028
rect 25044 17060 25096 17066
rect 25044 17002 25096 17008
rect 25056 16794 25084 17002
rect 25044 16788 25096 16794
rect 25044 16730 25096 16736
rect 25056 16182 25084 16730
rect 25044 16176 25096 16182
rect 25044 16118 25096 16124
rect 25044 15360 25096 15366
rect 25044 15302 25096 15308
rect 24952 13388 25004 13394
rect 24952 13330 25004 13336
rect 25056 13326 25084 15302
rect 24400 13320 24452 13326
rect 24400 13262 24452 13268
rect 25044 13320 25096 13326
rect 25044 13262 25096 13268
rect 25136 12844 25188 12850
rect 25136 12786 25188 12792
rect 25148 12238 25176 12786
rect 25136 12232 25188 12238
rect 25136 12174 25188 12180
rect 24860 12164 24912 12170
rect 24860 12106 24912 12112
rect 24872 11898 24900 12106
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 24400 11280 24452 11286
rect 24400 11222 24452 11228
rect 24412 6746 24440 11222
rect 24964 10470 24992 11698
rect 25148 11694 25176 12174
rect 25240 11898 25268 18566
rect 25228 11892 25280 11898
rect 25228 11834 25280 11840
rect 25136 11688 25188 11694
rect 25136 11630 25188 11636
rect 25516 11354 25544 22066
rect 25596 21344 25648 21350
rect 25596 21286 25648 21292
rect 25608 18358 25636 21286
rect 25700 20913 25728 23140
rect 25780 23044 25832 23050
rect 25780 22986 25832 22992
rect 25792 22166 25820 22986
rect 25780 22160 25832 22166
rect 25780 22102 25832 22108
rect 25780 21888 25832 21894
rect 25780 21830 25832 21836
rect 25686 20904 25742 20913
rect 25792 20874 25820 21830
rect 25686 20839 25742 20848
rect 25780 20868 25832 20874
rect 25700 20806 25728 20839
rect 25780 20810 25832 20816
rect 25688 20800 25740 20806
rect 25688 20742 25740 20748
rect 25596 18352 25648 18358
rect 25596 18294 25648 18300
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 25608 16998 25636 17138
rect 25596 16992 25648 16998
rect 25596 16934 25648 16940
rect 25608 15026 25636 16934
rect 25596 15020 25648 15026
rect 25596 14962 25648 14968
rect 25596 14000 25648 14006
rect 25596 13942 25648 13948
rect 25608 12238 25636 13942
rect 25688 13184 25740 13190
rect 25688 13126 25740 13132
rect 25700 12238 25728 13126
rect 25596 12232 25648 12238
rect 25596 12174 25648 12180
rect 25688 12232 25740 12238
rect 25688 12174 25740 12180
rect 25504 11348 25556 11354
rect 25504 11290 25556 11296
rect 25320 10668 25372 10674
rect 25320 10610 25372 10616
rect 25332 10470 25360 10610
rect 25516 10606 25544 11290
rect 25608 11150 25636 12174
rect 25688 11552 25740 11558
rect 25688 11494 25740 11500
rect 25596 11144 25648 11150
rect 25596 11086 25648 11092
rect 25700 11082 25728 11494
rect 25688 11076 25740 11082
rect 25688 11018 25740 11024
rect 25504 10600 25556 10606
rect 25504 10542 25556 10548
rect 24952 10464 25004 10470
rect 24952 10406 25004 10412
rect 25320 10464 25372 10470
rect 25320 10406 25372 10412
rect 25596 10464 25648 10470
rect 25596 10406 25648 10412
rect 25332 9722 25360 10406
rect 25320 9716 25372 9722
rect 25320 9658 25372 9664
rect 24952 9580 25004 9586
rect 24952 9522 25004 9528
rect 24504 8894 24900 8922
rect 24504 8498 24532 8894
rect 24872 8838 24900 8894
rect 24768 8832 24820 8838
rect 24768 8774 24820 8780
rect 24860 8832 24912 8838
rect 24860 8774 24912 8780
rect 24676 8560 24728 8566
rect 24676 8502 24728 8508
rect 24492 8492 24544 8498
rect 24492 8434 24544 8440
rect 24688 6934 24716 8502
rect 24780 8498 24808 8774
rect 24964 8634 24992 9522
rect 25412 9512 25464 9518
rect 25412 9454 25464 9460
rect 25228 9376 25280 9382
rect 25228 9318 25280 9324
rect 25136 8900 25188 8906
rect 25136 8842 25188 8848
rect 24952 8628 25004 8634
rect 24952 8570 25004 8576
rect 24768 8492 24820 8498
rect 24768 8434 24820 8440
rect 25044 8288 25096 8294
rect 25044 8230 25096 8236
rect 24860 7472 24912 7478
rect 24860 7414 24912 7420
rect 24676 6928 24728 6934
rect 24676 6870 24728 6876
rect 24676 6792 24728 6798
rect 24412 6730 24532 6746
rect 24676 6734 24728 6740
rect 24412 6724 24544 6730
rect 24412 6718 24492 6724
rect 24492 6666 24544 6672
rect 24688 6254 24716 6734
rect 24872 6390 24900 7414
rect 24952 7336 25004 7342
rect 24952 7278 25004 7284
rect 24964 6905 24992 7278
rect 24950 6896 25006 6905
rect 24950 6831 25006 6840
rect 24860 6384 24912 6390
rect 24860 6326 24912 6332
rect 24676 6248 24728 6254
rect 24676 6190 24728 6196
rect 24768 5840 24820 5846
rect 24768 5782 24820 5788
rect 24780 5710 24808 5782
rect 24872 5778 24900 6326
rect 24860 5772 24912 5778
rect 24860 5714 24912 5720
rect 24400 5704 24452 5710
rect 24400 5646 24452 5652
rect 24768 5704 24820 5710
rect 24768 5646 24820 5652
rect 24412 4826 24440 5646
rect 24492 5568 24544 5574
rect 24492 5510 24544 5516
rect 24504 5234 24532 5510
rect 24492 5228 24544 5234
rect 24492 5170 24544 5176
rect 24584 5024 24636 5030
rect 24584 4966 24636 4972
rect 24400 4820 24452 4826
rect 24400 4762 24452 4768
rect 24596 4690 24624 4966
rect 24584 4684 24636 4690
rect 24584 4626 24636 4632
rect 24400 4276 24452 4282
rect 24400 4218 24452 4224
rect 24412 3534 24440 4218
rect 24492 4140 24544 4146
rect 24492 4082 24544 4088
rect 24400 3528 24452 3534
rect 24400 3470 24452 3476
rect 24308 2576 24360 2582
rect 24308 2518 24360 2524
rect 24504 2514 24532 4082
rect 24596 3738 24624 4626
rect 24780 4214 24808 5646
rect 24768 4208 24820 4214
rect 24768 4150 24820 4156
rect 24964 4010 24992 6831
rect 25056 6662 25084 8230
rect 25148 8090 25176 8842
rect 25136 8084 25188 8090
rect 25136 8026 25188 8032
rect 25240 7886 25268 9318
rect 25424 9042 25452 9454
rect 25412 9036 25464 9042
rect 25412 8978 25464 8984
rect 25320 8900 25372 8906
rect 25320 8842 25372 8848
rect 25228 7880 25280 7886
rect 25228 7822 25280 7828
rect 25332 7750 25360 8842
rect 25608 8634 25636 10406
rect 25884 10266 25912 23598
rect 26068 22030 26096 23802
rect 26160 23730 26188 24074
rect 26148 23724 26200 23730
rect 26148 23666 26200 23672
rect 26252 23322 26280 25978
rect 26436 25974 26464 27406
rect 26516 27396 26568 27402
rect 26516 27338 26568 27344
rect 26528 26926 26556 27338
rect 26804 26994 26832 27610
rect 26792 26988 26844 26994
rect 26792 26930 26844 26936
rect 26976 26988 27028 26994
rect 26976 26930 27028 26936
rect 26516 26920 26568 26926
rect 26516 26862 26568 26868
rect 26424 25968 26476 25974
rect 26424 25910 26476 25916
rect 26884 25900 26936 25906
rect 26884 25842 26936 25848
rect 26424 25832 26476 25838
rect 26424 25774 26476 25780
rect 26332 25696 26384 25702
rect 26332 25638 26384 25644
rect 26240 23316 26292 23322
rect 26240 23258 26292 23264
rect 26056 22024 26108 22030
rect 26056 21966 26108 21972
rect 26148 22024 26200 22030
rect 26148 21966 26200 21972
rect 26160 21865 26188 21966
rect 26146 21856 26202 21865
rect 26146 21791 26202 21800
rect 26148 17536 26200 17542
rect 26148 17478 26200 17484
rect 26160 17202 26188 17478
rect 26148 17196 26200 17202
rect 26148 17138 26200 17144
rect 26344 17134 26372 25638
rect 26436 25294 26464 25774
rect 26792 25764 26844 25770
rect 26792 25706 26844 25712
rect 26804 25430 26832 25706
rect 26792 25424 26844 25430
rect 26792 25366 26844 25372
rect 26424 25288 26476 25294
rect 26424 25230 26476 25236
rect 26700 25288 26752 25294
rect 26700 25230 26752 25236
rect 26436 24750 26464 25230
rect 26712 24954 26740 25230
rect 26804 25226 26832 25366
rect 26792 25220 26844 25226
rect 26792 25162 26844 25168
rect 26700 24948 26752 24954
rect 26700 24890 26752 24896
rect 26608 24880 26660 24886
rect 26608 24822 26660 24828
rect 26424 24744 26476 24750
rect 26424 24686 26476 24692
rect 26516 24676 26568 24682
rect 26516 24618 26568 24624
rect 26424 23724 26476 23730
rect 26424 23666 26476 23672
rect 26436 23118 26464 23666
rect 26424 23112 26476 23118
rect 26424 23054 26476 23060
rect 26436 22778 26464 23054
rect 26424 22772 26476 22778
rect 26424 22714 26476 22720
rect 26436 22166 26464 22714
rect 26424 22160 26476 22166
rect 26424 22102 26476 22108
rect 26528 22098 26556 24618
rect 26516 22092 26568 22098
rect 26516 22034 26568 22040
rect 26528 20942 26556 22034
rect 26620 22030 26648 24822
rect 26792 24812 26844 24818
rect 26792 24754 26844 24760
rect 26804 24206 26832 24754
rect 26896 24682 26924 25842
rect 26988 25158 27016 26930
rect 27068 25900 27120 25906
rect 27068 25842 27120 25848
rect 27080 25498 27108 25842
rect 27068 25492 27120 25498
rect 27068 25434 27120 25440
rect 26976 25152 27028 25158
rect 26976 25094 27028 25100
rect 26884 24676 26936 24682
rect 26884 24618 26936 24624
rect 26896 24342 26924 24618
rect 26884 24336 26936 24342
rect 26884 24278 26936 24284
rect 26792 24200 26844 24206
rect 26792 24142 26844 24148
rect 26700 24132 26752 24138
rect 26700 24074 26752 24080
rect 26712 23798 26740 24074
rect 26700 23792 26752 23798
rect 26700 23734 26752 23740
rect 26608 22024 26660 22030
rect 26608 21966 26660 21972
rect 26516 20936 26568 20942
rect 26516 20878 26568 20884
rect 26608 20800 26660 20806
rect 26608 20742 26660 20748
rect 26516 20256 26568 20262
rect 26516 20198 26568 20204
rect 26332 17128 26384 17134
rect 26332 17070 26384 17076
rect 26148 17060 26200 17066
rect 26148 17002 26200 17008
rect 26160 16590 26188 17002
rect 26148 16584 26200 16590
rect 26148 16526 26200 16532
rect 26148 16108 26200 16114
rect 26148 16050 26200 16056
rect 26160 15706 26188 16050
rect 26148 15700 26200 15706
rect 26148 15642 26200 15648
rect 26148 15496 26200 15502
rect 26148 15438 26200 15444
rect 26160 15026 26188 15438
rect 26148 15020 26200 15026
rect 26148 14962 26200 14968
rect 26160 14482 26188 14962
rect 26148 14476 26200 14482
rect 26148 14418 26200 14424
rect 26056 13728 26108 13734
rect 26056 13670 26108 13676
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 26068 13462 26096 13670
rect 26056 13456 26108 13462
rect 26056 13398 26108 13404
rect 26252 13326 26280 13670
rect 26424 13524 26476 13530
rect 26424 13466 26476 13472
rect 26240 13320 26292 13326
rect 26240 13262 26292 13268
rect 26436 12170 26464 13466
rect 26528 13394 26556 20198
rect 26620 18766 26648 20742
rect 26700 20392 26752 20398
rect 26700 20334 26752 20340
rect 26712 19854 26740 20334
rect 26700 19848 26752 19854
rect 26700 19790 26752 19796
rect 26700 19712 26752 19718
rect 26700 19654 26752 19660
rect 26712 19446 26740 19654
rect 26700 19440 26752 19446
rect 26700 19382 26752 19388
rect 26608 18760 26660 18766
rect 26608 18702 26660 18708
rect 26620 17218 26648 18702
rect 26620 17190 26740 17218
rect 26608 14816 26660 14822
rect 26608 14758 26660 14764
rect 26516 13388 26568 13394
rect 26516 13330 26568 13336
rect 26424 12164 26476 12170
rect 26424 12106 26476 12112
rect 25964 12096 26016 12102
rect 25964 12038 26016 12044
rect 25872 10260 25924 10266
rect 25872 10202 25924 10208
rect 25884 9654 25912 10202
rect 25872 9648 25924 9654
rect 25872 9590 25924 9596
rect 25596 8628 25648 8634
rect 25596 8570 25648 8576
rect 25412 8492 25464 8498
rect 25412 8434 25464 8440
rect 25320 7744 25372 7750
rect 25320 7686 25372 7692
rect 25424 7478 25452 8434
rect 25412 7472 25464 7478
rect 25412 7414 25464 7420
rect 25136 7336 25188 7342
rect 25136 7278 25188 7284
rect 25148 7002 25176 7278
rect 25320 7200 25372 7206
rect 25320 7142 25372 7148
rect 25136 6996 25188 7002
rect 25136 6938 25188 6944
rect 25044 6656 25096 6662
rect 25044 6598 25096 6604
rect 25332 6322 25360 7142
rect 25044 6316 25096 6322
rect 25044 6258 25096 6264
rect 25320 6316 25372 6322
rect 25320 6258 25372 6264
rect 25056 5302 25084 6258
rect 25136 5840 25188 5846
rect 25136 5782 25188 5788
rect 25044 5296 25096 5302
rect 25044 5238 25096 5244
rect 24860 4004 24912 4010
rect 24860 3946 24912 3952
rect 24952 4004 25004 4010
rect 24952 3946 25004 3952
rect 24584 3732 24636 3738
rect 24584 3674 24636 3680
rect 24872 3058 24900 3946
rect 24964 3602 24992 3946
rect 24952 3596 25004 3602
rect 24952 3538 25004 3544
rect 24952 3188 25004 3194
rect 24952 3130 25004 3136
rect 24860 3052 24912 3058
rect 24860 2994 24912 3000
rect 24964 2938 24992 3130
rect 25056 3058 25084 5238
rect 25044 3052 25096 3058
rect 25044 2994 25096 3000
rect 24872 2910 24992 2938
rect 24492 2508 24544 2514
rect 24492 2450 24544 2456
rect 24872 2378 24900 2910
rect 25148 2774 25176 5782
rect 25412 5024 25464 5030
rect 25412 4966 25464 4972
rect 25424 4826 25452 4966
rect 25412 4820 25464 4826
rect 25412 4762 25464 4768
rect 25596 4616 25648 4622
rect 25596 4558 25648 4564
rect 25320 4480 25372 4486
rect 25320 4422 25372 4428
rect 25228 3528 25280 3534
rect 25228 3470 25280 3476
rect 25240 3194 25268 3470
rect 25228 3188 25280 3194
rect 25228 3130 25280 3136
rect 24964 2746 25176 2774
rect 24860 2372 24912 2378
rect 24860 2314 24912 2320
rect 24216 2304 24268 2310
rect 24216 2246 24268 2252
rect 24228 800 24256 2246
rect 24584 1420 24636 1426
rect 24584 1362 24636 1368
rect 24596 800 24624 1362
rect 24964 800 24992 2746
rect 25240 2446 25268 3130
rect 25332 3058 25360 4422
rect 25412 3936 25464 3942
rect 25412 3878 25464 3884
rect 25320 3052 25372 3058
rect 25320 2994 25372 3000
rect 25424 2774 25452 3878
rect 25332 2746 25452 2774
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 25332 800 25360 2746
rect 25608 2650 25636 4558
rect 25976 4146 26004 12038
rect 26240 11144 26292 11150
rect 26240 11086 26292 11092
rect 26252 10062 26280 11086
rect 26240 10056 26292 10062
rect 26240 9998 26292 10004
rect 26148 9988 26200 9994
rect 26148 9930 26200 9936
rect 26160 9722 26188 9930
rect 26148 9716 26200 9722
rect 26148 9658 26200 9664
rect 26252 9625 26280 9998
rect 26332 9920 26384 9926
rect 26332 9862 26384 9868
rect 26238 9616 26294 9625
rect 26344 9586 26372 9862
rect 26238 9551 26294 9560
rect 26332 9580 26384 9586
rect 26252 8974 26280 9551
rect 26620 9568 26648 14758
rect 26712 12434 26740 17190
rect 26804 13818 26832 24142
rect 26988 21078 27016 25094
rect 27068 24812 27120 24818
rect 27068 24754 27120 24760
rect 27080 24410 27108 24754
rect 27068 24404 27120 24410
rect 27068 24346 27120 24352
rect 27172 23594 27200 27662
rect 27528 27600 27580 27606
rect 27528 27542 27580 27548
rect 27252 27328 27304 27334
rect 27252 27270 27304 27276
rect 27264 27062 27292 27270
rect 27252 27056 27304 27062
rect 27252 26998 27304 27004
rect 27160 23588 27212 23594
rect 27160 23530 27212 23536
rect 27344 22568 27396 22574
rect 27344 22510 27396 22516
rect 27160 21548 27212 21554
rect 27212 21508 27292 21536
rect 27160 21490 27212 21496
rect 27068 21344 27120 21350
rect 27068 21286 27120 21292
rect 26976 21072 27028 21078
rect 26976 21014 27028 21020
rect 27080 20874 27108 21286
rect 27068 20868 27120 20874
rect 27068 20810 27120 20816
rect 26884 20596 26936 20602
rect 26884 20538 26936 20544
rect 26896 19854 26924 20538
rect 27264 20534 27292 21508
rect 27252 20528 27304 20534
rect 27252 20470 27304 20476
rect 26976 20256 27028 20262
rect 26976 20198 27028 20204
rect 26884 19848 26936 19854
rect 26884 19790 26936 19796
rect 26988 18766 27016 20198
rect 27160 19712 27212 19718
rect 27160 19654 27212 19660
rect 27068 19372 27120 19378
rect 27068 19314 27120 19320
rect 27080 18970 27108 19314
rect 27068 18964 27120 18970
rect 27068 18906 27120 18912
rect 26976 18760 27028 18766
rect 26976 18702 27028 18708
rect 26976 17604 27028 17610
rect 26976 17546 27028 17552
rect 26988 17338 27016 17546
rect 26976 17332 27028 17338
rect 26976 17274 27028 17280
rect 27068 16652 27120 16658
rect 27068 16594 27120 16600
rect 27080 16114 27108 16594
rect 27172 16538 27200 19654
rect 27264 18766 27292 20470
rect 27356 19825 27384 22510
rect 27436 21548 27488 21554
rect 27436 21490 27488 21496
rect 27448 20505 27476 21490
rect 27434 20496 27490 20505
rect 27434 20431 27490 20440
rect 27448 19854 27476 20431
rect 27436 19848 27488 19854
rect 27342 19816 27398 19825
rect 27436 19790 27488 19796
rect 27342 19751 27398 19760
rect 27356 18902 27384 19751
rect 27436 19712 27488 19718
rect 27436 19654 27488 19660
rect 27448 19446 27476 19654
rect 27436 19440 27488 19446
rect 27436 19382 27488 19388
rect 27344 18896 27396 18902
rect 27344 18838 27396 18844
rect 27252 18760 27304 18766
rect 27252 18702 27304 18708
rect 27264 18290 27292 18702
rect 27252 18284 27304 18290
rect 27252 18226 27304 18232
rect 27252 17128 27304 17134
rect 27252 17070 27304 17076
rect 27264 16658 27292 17070
rect 27252 16652 27304 16658
rect 27252 16594 27304 16600
rect 27172 16510 27292 16538
rect 27068 16108 27120 16114
rect 27068 16050 27120 16056
rect 26976 15360 27028 15366
rect 26976 15302 27028 15308
rect 26988 14414 27016 15302
rect 26976 14408 27028 14414
rect 26976 14350 27028 14356
rect 27160 14408 27212 14414
rect 27160 14350 27212 14356
rect 27068 14272 27120 14278
rect 27068 14214 27120 14220
rect 27080 13938 27108 14214
rect 27068 13932 27120 13938
rect 27068 13874 27120 13880
rect 26804 13790 27108 13818
rect 26976 13320 27028 13326
rect 26976 13262 27028 13268
rect 26884 13252 26936 13258
rect 26884 13194 26936 13200
rect 26712 12406 26832 12434
rect 26700 10464 26752 10470
rect 26700 10406 26752 10412
rect 26712 10198 26740 10406
rect 26700 10192 26752 10198
rect 26700 10134 26752 10140
rect 26620 9540 26740 9568
rect 26332 9522 26384 9528
rect 26608 9444 26660 9450
rect 26608 9386 26660 9392
rect 26240 8968 26292 8974
rect 26240 8910 26292 8916
rect 26516 8832 26568 8838
rect 26516 8774 26568 8780
rect 26424 8492 26476 8498
rect 26424 8434 26476 8440
rect 26240 7948 26292 7954
rect 26240 7890 26292 7896
rect 26252 6798 26280 7890
rect 26436 7478 26464 8434
rect 26424 7472 26476 7478
rect 26424 7414 26476 7420
rect 26332 7404 26384 7410
rect 26332 7346 26384 7352
rect 26240 6792 26292 6798
rect 26240 6734 26292 6740
rect 26056 6724 26108 6730
rect 26056 6666 26108 6672
rect 25964 4140 26016 4146
rect 25964 4082 26016 4088
rect 25688 4072 25740 4078
rect 25688 4014 25740 4020
rect 25596 2644 25648 2650
rect 25596 2586 25648 2592
rect 25504 2372 25556 2378
rect 25504 2314 25556 2320
rect 25516 2106 25544 2314
rect 25504 2100 25556 2106
rect 25504 2042 25556 2048
rect 25700 800 25728 4014
rect 25780 2848 25832 2854
rect 25780 2790 25832 2796
rect 25792 2446 25820 2790
rect 25780 2440 25832 2446
rect 25780 2382 25832 2388
rect 25792 1970 25820 2382
rect 25780 1964 25832 1970
rect 25780 1906 25832 1912
rect 26068 800 26096 6666
rect 26240 6452 26292 6458
rect 26240 6394 26292 6400
rect 26252 5574 26280 6394
rect 26344 5914 26372 7346
rect 26424 6996 26476 7002
rect 26528 6984 26556 8774
rect 26476 6956 26556 6984
rect 26424 6938 26476 6944
rect 26332 5908 26384 5914
rect 26332 5850 26384 5856
rect 26436 5794 26464 6938
rect 26516 6112 26568 6118
rect 26516 6054 26568 6060
rect 26344 5766 26464 5794
rect 26344 5710 26372 5766
rect 26528 5710 26556 6054
rect 26332 5704 26384 5710
rect 26332 5646 26384 5652
rect 26516 5704 26568 5710
rect 26516 5646 26568 5652
rect 26424 5636 26476 5642
rect 26424 5578 26476 5584
rect 26240 5568 26292 5574
rect 26240 5510 26292 5516
rect 26252 5386 26280 5510
rect 26252 5358 26372 5386
rect 26240 5228 26292 5234
rect 26240 5170 26292 5176
rect 26252 4826 26280 5170
rect 26240 4820 26292 4826
rect 26240 4762 26292 4768
rect 26344 4690 26372 5358
rect 26436 5234 26464 5578
rect 26424 5228 26476 5234
rect 26424 5170 26476 5176
rect 26332 4684 26384 4690
rect 26332 4626 26384 4632
rect 26240 4208 26292 4214
rect 26240 4150 26292 4156
rect 26252 3738 26280 4150
rect 26424 3936 26476 3942
rect 26424 3878 26476 3884
rect 26240 3732 26292 3738
rect 26240 3674 26292 3680
rect 26436 800 26464 3878
rect 26620 2038 26648 9386
rect 26712 3534 26740 9540
rect 26804 8294 26832 12406
rect 26896 11762 26924 13194
rect 26988 12442 27016 13262
rect 26976 12436 27028 12442
rect 26976 12378 27028 12384
rect 26884 11756 26936 11762
rect 26884 11698 26936 11704
rect 26976 10532 27028 10538
rect 26976 10474 27028 10480
rect 26988 9586 27016 10474
rect 26976 9580 27028 9586
rect 26976 9522 27028 9528
rect 26884 9036 26936 9042
rect 26884 8978 26936 8984
rect 26896 8412 26924 8978
rect 26896 8384 27016 8412
rect 26792 8288 26844 8294
rect 26792 8230 26844 8236
rect 26804 7954 26832 8230
rect 26792 7948 26844 7954
rect 26792 7890 26844 7896
rect 26884 7880 26936 7886
rect 26884 7822 26936 7828
rect 26896 7410 26924 7822
rect 26884 7404 26936 7410
rect 26884 7346 26936 7352
rect 26896 5846 26924 7346
rect 26988 7342 27016 8384
rect 26976 7336 27028 7342
rect 26976 7278 27028 7284
rect 26976 6996 27028 7002
rect 26976 6938 27028 6944
rect 26988 6390 27016 6938
rect 27080 6458 27108 13790
rect 27172 13530 27200 14350
rect 27160 13524 27212 13530
rect 27160 13466 27212 13472
rect 27264 13394 27292 16510
rect 27540 16182 27568 27542
rect 27632 25974 27660 27814
rect 27896 27600 27948 27606
rect 27896 27542 27948 27548
rect 27804 27464 27856 27470
rect 27804 27406 27856 27412
rect 27712 27396 27764 27402
rect 27712 27338 27764 27344
rect 27724 27062 27752 27338
rect 27816 27305 27844 27406
rect 27802 27296 27858 27305
rect 27802 27231 27858 27240
rect 27712 27056 27764 27062
rect 27712 26998 27764 27004
rect 27724 26382 27752 26998
rect 27908 26994 27936 27542
rect 27896 26988 27948 26994
rect 27896 26930 27948 26936
rect 27804 26920 27856 26926
rect 27804 26862 27856 26868
rect 27712 26376 27764 26382
rect 27712 26318 27764 26324
rect 27620 25968 27672 25974
rect 27620 25910 27672 25916
rect 27712 25288 27764 25294
rect 27710 25256 27712 25265
rect 27764 25256 27766 25265
rect 27710 25191 27766 25200
rect 27712 23520 27764 23526
rect 27712 23462 27764 23468
rect 27724 22522 27752 23462
rect 27632 22494 27752 22522
rect 27632 17218 27660 22494
rect 27712 22432 27764 22438
rect 27712 22374 27764 22380
rect 27724 21962 27752 22374
rect 27692 21956 27752 21962
rect 27744 21916 27752 21956
rect 27692 21898 27744 21904
rect 27710 21720 27766 21729
rect 27710 21655 27712 21664
rect 27764 21655 27766 21664
rect 27712 21626 27764 21632
rect 27710 21584 27766 21593
rect 27710 21519 27766 21528
rect 27724 21078 27752 21519
rect 27712 21072 27764 21078
rect 27712 21014 27764 21020
rect 27816 20602 27844 26862
rect 27896 25288 27948 25294
rect 27896 25230 27948 25236
rect 27908 24954 27936 25230
rect 27896 24948 27948 24954
rect 27896 24890 27948 24896
rect 27908 23730 27936 24890
rect 27896 23724 27948 23730
rect 27896 23666 27948 23672
rect 27896 22636 27948 22642
rect 27896 22578 27948 22584
rect 27908 21729 27936 22578
rect 27894 21720 27950 21729
rect 27894 21655 27950 21664
rect 27894 21584 27950 21593
rect 27894 21519 27896 21528
rect 27948 21519 27950 21528
rect 27896 21490 27948 21496
rect 27804 20596 27856 20602
rect 27804 20538 27856 20544
rect 27804 20460 27856 20466
rect 27804 20402 27856 20408
rect 27712 19984 27764 19990
rect 27712 19926 27764 19932
rect 27724 17728 27752 19926
rect 27816 19514 27844 20402
rect 27896 19848 27948 19854
rect 27896 19790 27948 19796
rect 27804 19508 27856 19514
rect 27804 19450 27856 19456
rect 27908 18970 27936 19790
rect 27896 18964 27948 18970
rect 27896 18906 27948 18912
rect 27724 17700 27936 17728
rect 27632 17190 27844 17218
rect 27620 16516 27672 16522
rect 27620 16458 27672 16464
rect 27528 16176 27580 16182
rect 27528 16118 27580 16124
rect 27632 15706 27660 16458
rect 27712 15904 27764 15910
rect 27712 15846 27764 15852
rect 27620 15700 27672 15706
rect 27620 15642 27672 15648
rect 27724 15586 27752 15846
rect 27632 15558 27752 15586
rect 27528 15496 27580 15502
rect 27632 15484 27660 15558
rect 27580 15456 27660 15484
rect 27528 15438 27580 15444
rect 27528 14340 27580 14346
rect 27528 14282 27580 14288
rect 27252 13388 27304 13394
rect 27252 13330 27304 13336
rect 27540 13326 27568 14282
rect 27528 13320 27580 13326
rect 27528 13262 27580 13268
rect 27632 11830 27660 15456
rect 27712 13932 27764 13938
rect 27712 13874 27764 13880
rect 27724 13530 27752 13874
rect 27712 13524 27764 13530
rect 27712 13466 27764 13472
rect 27816 12434 27844 17190
rect 27908 17116 27936 17700
rect 28000 17218 28028 28358
rect 28080 27396 28132 27402
rect 28080 27338 28132 27344
rect 28092 26858 28120 27338
rect 28184 26926 28212 32422
rect 28356 32370 28408 32376
rect 28368 31482 28396 32370
rect 28356 31476 28408 31482
rect 28356 31418 28408 31424
rect 28356 30796 28408 30802
rect 28356 30738 28408 30744
rect 28264 30048 28316 30054
rect 28264 29990 28316 29996
rect 28276 27606 28304 29990
rect 28368 29102 28396 30738
rect 28356 29096 28408 29102
rect 28356 29038 28408 29044
rect 28356 28484 28408 28490
rect 28356 28426 28408 28432
rect 28368 28082 28396 28426
rect 28356 28076 28408 28082
rect 28356 28018 28408 28024
rect 28264 27600 28316 27606
rect 28264 27542 28316 27548
rect 28264 27464 28316 27470
rect 28262 27432 28264 27441
rect 28316 27432 28318 27441
rect 28262 27367 28318 27376
rect 28172 26920 28224 26926
rect 28172 26862 28224 26868
rect 28080 26852 28132 26858
rect 28080 26794 28132 26800
rect 28092 23730 28120 26794
rect 28172 25696 28224 25702
rect 28172 25638 28224 25644
rect 28184 25294 28212 25638
rect 28172 25288 28224 25294
rect 28172 25230 28224 25236
rect 28276 24256 28304 27367
rect 28354 27296 28410 27305
rect 28354 27231 28410 27240
rect 28368 27062 28396 27231
rect 28356 27056 28408 27062
rect 28356 26998 28408 27004
rect 28460 24410 28488 35550
rect 28540 35556 28592 35562
rect 28540 35498 28592 35504
rect 28540 35080 28592 35086
rect 28540 35022 28592 35028
rect 28552 34610 28580 35022
rect 28540 34604 28592 34610
rect 28540 34546 28592 34552
rect 28552 33318 28580 34546
rect 28540 33312 28592 33318
rect 28540 33254 28592 33260
rect 28552 32298 28580 33254
rect 28736 33114 28764 35634
rect 28724 33108 28776 33114
rect 28724 33050 28776 33056
rect 28736 32570 28764 33050
rect 28724 32564 28776 32570
rect 28724 32506 28776 32512
rect 28540 32292 28592 32298
rect 28540 32234 28592 32240
rect 28552 27538 28580 32234
rect 28632 31136 28684 31142
rect 28632 31078 28684 31084
rect 28644 30734 28672 31078
rect 28632 30728 28684 30734
rect 28632 30670 28684 30676
rect 28540 27532 28592 27538
rect 28540 27474 28592 27480
rect 28644 27402 28672 30670
rect 28632 27396 28684 27402
rect 28632 27338 28684 27344
rect 28540 27328 28592 27334
rect 28540 27270 28592 27276
rect 28448 24404 28500 24410
rect 28448 24346 28500 24352
rect 28184 24228 28304 24256
rect 28080 23724 28132 23730
rect 28080 23666 28132 23672
rect 28184 23610 28212 24228
rect 28448 24200 28500 24206
rect 28448 24142 28500 24148
rect 28264 24132 28316 24138
rect 28264 24074 28316 24080
rect 28276 23866 28304 24074
rect 28356 24064 28408 24070
rect 28356 24006 28408 24012
rect 28264 23860 28316 23866
rect 28264 23802 28316 23808
rect 28264 23724 28316 23730
rect 28264 23666 28316 23672
rect 28092 23582 28212 23610
rect 28092 22545 28120 23582
rect 28078 22536 28134 22545
rect 28078 22471 28134 22480
rect 28080 22432 28132 22438
rect 28080 22374 28132 22380
rect 28092 21418 28120 22374
rect 28276 21690 28304 23666
rect 28368 22642 28396 24006
rect 28460 23526 28488 24142
rect 28448 23520 28500 23526
rect 28448 23462 28500 23468
rect 28460 23118 28488 23462
rect 28448 23112 28500 23118
rect 28448 23054 28500 23060
rect 28356 22636 28408 22642
rect 28356 22578 28408 22584
rect 28354 22536 28410 22545
rect 28354 22471 28410 22480
rect 28264 21684 28316 21690
rect 28264 21626 28316 21632
rect 28368 21554 28396 22471
rect 28448 22228 28500 22234
rect 28448 22170 28500 22176
rect 28460 21622 28488 22170
rect 28448 21616 28500 21622
rect 28448 21558 28500 21564
rect 28356 21548 28408 21554
rect 28356 21490 28408 21496
rect 28080 21412 28132 21418
rect 28080 21354 28132 21360
rect 28264 21344 28316 21350
rect 28264 21286 28316 21292
rect 28172 21004 28224 21010
rect 28172 20946 28224 20952
rect 28078 20904 28134 20913
rect 28078 20839 28080 20848
rect 28132 20839 28134 20848
rect 28080 20810 28132 20816
rect 28078 20632 28134 20641
rect 28078 20567 28134 20576
rect 28092 20466 28120 20567
rect 28080 20460 28132 20466
rect 28080 20402 28132 20408
rect 28092 18766 28120 20402
rect 28184 19990 28212 20946
rect 28172 19984 28224 19990
rect 28172 19926 28224 19932
rect 28172 19848 28224 19854
rect 28172 19790 28224 19796
rect 28184 18834 28212 19790
rect 28172 18828 28224 18834
rect 28172 18770 28224 18776
rect 28080 18760 28132 18766
rect 28080 18702 28132 18708
rect 28172 17740 28224 17746
rect 28172 17682 28224 17688
rect 28000 17190 28120 17218
rect 27908 17088 28028 17116
rect 27896 15972 27948 15978
rect 27896 15914 27948 15920
rect 27908 14618 27936 15914
rect 27896 14612 27948 14618
rect 27896 14554 27948 14560
rect 28000 14498 28028 17088
rect 27724 12406 27844 12434
rect 27908 14470 28028 14498
rect 27620 11824 27672 11830
rect 27620 11766 27672 11772
rect 27344 11552 27396 11558
rect 27344 11494 27396 11500
rect 27252 9376 27304 9382
rect 27252 9318 27304 9324
rect 27264 8906 27292 9318
rect 27252 8900 27304 8906
rect 27252 8842 27304 8848
rect 27252 7744 27304 7750
rect 27252 7686 27304 7692
rect 27264 7410 27292 7686
rect 27252 7404 27304 7410
rect 27252 7346 27304 7352
rect 27068 6452 27120 6458
rect 27068 6394 27120 6400
rect 26976 6384 27028 6390
rect 26976 6326 27028 6332
rect 26884 5840 26936 5846
rect 26884 5782 26936 5788
rect 26884 5704 26936 5710
rect 26884 5646 26936 5652
rect 26792 5568 26844 5574
rect 26792 5510 26844 5516
rect 26804 4622 26832 5510
rect 26792 4616 26844 4622
rect 26792 4558 26844 4564
rect 26700 3528 26752 3534
rect 26700 3470 26752 3476
rect 26608 2032 26660 2038
rect 26608 1974 26660 1980
rect 26896 800 26924 5646
rect 26988 5166 27016 6326
rect 27080 6322 27108 6394
rect 27068 6316 27120 6322
rect 27068 6258 27120 6264
rect 26976 5160 27028 5166
rect 26976 5102 27028 5108
rect 27356 4146 27384 11494
rect 27528 11076 27580 11082
rect 27528 11018 27580 11024
rect 27436 10464 27488 10470
rect 27436 10406 27488 10412
rect 27448 10062 27476 10406
rect 27540 10266 27568 11018
rect 27620 10804 27672 10810
rect 27620 10746 27672 10752
rect 27528 10260 27580 10266
rect 27528 10202 27580 10208
rect 27436 10056 27488 10062
rect 27436 9998 27488 10004
rect 27526 9616 27582 9625
rect 27526 9551 27582 9560
rect 27540 9518 27568 9551
rect 27528 9512 27580 9518
rect 27528 9454 27580 9460
rect 27540 8566 27568 9454
rect 27528 8560 27580 8566
rect 27528 8502 27580 8508
rect 27540 7886 27568 8502
rect 27528 7880 27580 7886
rect 27528 7822 27580 7828
rect 27540 7002 27568 7822
rect 27528 6996 27580 7002
rect 27528 6938 27580 6944
rect 27632 6730 27660 10746
rect 27724 8566 27752 12406
rect 27804 12232 27856 12238
rect 27804 12174 27856 12180
rect 27816 11694 27844 12174
rect 27804 11688 27856 11694
rect 27804 11630 27856 11636
rect 27908 11354 27936 14470
rect 27988 14408 28040 14414
rect 27988 14350 28040 14356
rect 28000 13938 28028 14350
rect 27988 13932 28040 13938
rect 27988 13874 28040 13880
rect 27896 11348 27948 11354
rect 27896 11290 27948 11296
rect 27908 10826 27936 11290
rect 27816 10798 27936 10826
rect 27816 10742 27844 10798
rect 27804 10736 27856 10742
rect 27804 10678 27856 10684
rect 27804 8832 27856 8838
rect 27804 8774 27856 8780
rect 27988 8832 28040 8838
rect 27988 8774 28040 8780
rect 27712 8560 27764 8566
rect 27712 8502 27764 8508
rect 27816 8498 27844 8774
rect 27804 8492 27856 8498
rect 27804 8434 27856 8440
rect 27804 7812 27856 7818
rect 27804 7754 27856 7760
rect 27712 7744 27764 7750
rect 27712 7686 27764 7692
rect 27620 6724 27672 6730
rect 27620 6666 27672 6672
rect 27436 6316 27488 6322
rect 27436 6258 27488 6264
rect 27620 6316 27672 6322
rect 27620 6258 27672 6264
rect 27448 5778 27476 6258
rect 27632 5914 27660 6258
rect 27620 5908 27672 5914
rect 27620 5850 27672 5856
rect 27436 5772 27488 5778
rect 27436 5714 27488 5720
rect 27724 5710 27752 7686
rect 27816 7206 27844 7754
rect 28000 7410 28028 8774
rect 28092 7818 28120 17190
rect 28184 16046 28212 17682
rect 28172 16040 28224 16046
rect 28172 15982 28224 15988
rect 28172 15904 28224 15910
rect 28172 15846 28224 15852
rect 28184 15502 28212 15846
rect 28172 15496 28224 15502
rect 28172 15438 28224 15444
rect 28276 14482 28304 21286
rect 28368 20534 28396 21490
rect 28448 20800 28500 20806
rect 28448 20742 28500 20748
rect 28356 20528 28408 20534
rect 28460 20505 28488 20742
rect 28356 20470 28408 20476
rect 28446 20496 28502 20505
rect 28446 20431 28502 20440
rect 28448 19916 28500 19922
rect 28448 19858 28500 19864
rect 28354 19816 28410 19825
rect 28354 19751 28356 19760
rect 28408 19751 28410 19760
rect 28356 19722 28408 19728
rect 28460 19689 28488 19858
rect 28446 19680 28502 19689
rect 28446 19615 28502 19624
rect 28356 17672 28408 17678
rect 28356 17614 28408 17620
rect 28368 17338 28396 17614
rect 28356 17332 28408 17338
rect 28356 17274 28408 17280
rect 28356 16448 28408 16454
rect 28356 16390 28408 16396
rect 28368 16114 28396 16390
rect 28356 16108 28408 16114
rect 28356 16050 28408 16056
rect 28448 16108 28500 16114
rect 28448 16050 28500 16056
rect 28460 15026 28488 16050
rect 28552 16046 28580 27270
rect 28736 26994 28764 32506
rect 28828 31754 28856 35634
rect 28920 34610 28948 37266
rect 29564 36582 29592 37606
rect 29840 36922 29868 46990
rect 30392 46918 30420 49200
rect 30748 47456 30800 47462
rect 30748 47398 30800 47404
rect 30760 47258 30788 47398
rect 30748 47252 30800 47258
rect 30748 47194 30800 47200
rect 31024 47184 31076 47190
rect 31024 47126 31076 47132
rect 30380 46912 30432 46918
rect 30380 46854 30432 46860
rect 29920 46504 29972 46510
rect 29920 46446 29972 46452
rect 29828 36916 29880 36922
rect 29828 36858 29880 36864
rect 29552 36576 29604 36582
rect 29552 36518 29604 36524
rect 29932 36310 29960 46446
rect 30380 45484 30432 45490
rect 30380 45426 30432 45432
rect 29920 36304 29972 36310
rect 29920 36246 29972 36252
rect 29736 35692 29788 35698
rect 29736 35634 29788 35640
rect 29092 35080 29144 35086
rect 29092 35022 29144 35028
rect 28908 34604 28960 34610
rect 28908 34546 28960 34552
rect 29104 34542 29132 35022
rect 29748 34746 29776 35634
rect 30392 35290 30420 45426
rect 30564 35760 30616 35766
rect 30564 35702 30616 35708
rect 30380 35284 30432 35290
rect 30380 35226 30432 35232
rect 30196 35216 30248 35222
rect 30196 35158 30248 35164
rect 30472 35216 30524 35222
rect 30472 35158 30524 35164
rect 29736 34740 29788 34746
rect 29736 34682 29788 34688
rect 29092 34536 29144 34542
rect 29092 34478 29144 34484
rect 29000 33516 29052 33522
rect 29000 33458 29052 33464
rect 28828 31726 28948 31754
rect 28816 30388 28868 30394
rect 28816 30330 28868 30336
rect 28724 26988 28776 26994
rect 28724 26930 28776 26936
rect 28632 25152 28684 25158
rect 28632 25094 28684 25100
rect 28644 17746 28672 25094
rect 28724 24064 28776 24070
rect 28724 24006 28776 24012
rect 28736 23866 28764 24006
rect 28724 23860 28776 23866
rect 28724 23802 28776 23808
rect 28724 23724 28776 23730
rect 28724 23666 28776 23672
rect 28736 23322 28764 23666
rect 28724 23316 28776 23322
rect 28724 23258 28776 23264
rect 28828 22137 28856 30330
rect 28920 30054 28948 31726
rect 29012 31414 29040 33458
rect 29000 31408 29052 31414
rect 29000 31350 29052 31356
rect 28908 30048 28960 30054
rect 28908 29990 28960 29996
rect 28908 29844 28960 29850
rect 28908 29786 28960 29792
rect 28920 29034 28948 29786
rect 28908 29028 28960 29034
rect 28908 28970 28960 28976
rect 28920 27062 28948 28970
rect 29000 28416 29052 28422
rect 29000 28358 29052 28364
rect 29012 28218 29040 28358
rect 29000 28212 29052 28218
rect 29000 28154 29052 28160
rect 29000 28008 29052 28014
rect 29000 27950 29052 27956
rect 29012 27130 29040 27950
rect 29104 27130 29132 34478
rect 29644 34468 29696 34474
rect 29644 34410 29696 34416
rect 29552 33992 29604 33998
rect 29552 33934 29604 33940
rect 29564 33522 29592 33934
rect 29552 33516 29604 33522
rect 29552 33458 29604 33464
rect 29184 31340 29236 31346
rect 29184 31282 29236 31288
rect 29196 30326 29224 31282
rect 29184 30320 29236 30326
rect 29184 30262 29236 30268
rect 29564 29850 29592 33458
rect 29656 31958 29684 34410
rect 30208 34134 30236 35158
rect 30380 34944 30432 34950
rect 30380 34886 30432 34892
rect 30392 34626 30420 34886
rect 30300 34610 30420 34626
rect 30288 34604 30420 34610
rect 30340 34598 30420 34604
rect 30288 34546 30340 34552
rect 30196 34128 30248 34134
rect 30196 34070 30248 34076
rect 30288 33856 30340 33862
rect 30288 33798 30340 33804
rect 30300 33590 30328 33798
rect 30380 33652 30432 33658
rect 30380 33594 30432 33600
rect 30288 33584 30340 33590
rect 30288 33526 30340 33532
rect 30196 32360 30248 32366
rect 30196 32302 30248 32308
rect 29644 31952 29696 31958
rect 29644 31894 29696 31900
rect 30208 31754 30236 32302
rect 30116 31726 30236 31754
rect 30116 31414 30144 31726
rect 30104 31408 30156 31414
rect 30104 31350 30156 31356
rect 29552 29844 29604 29850
rect 29552 29786 29604 29792
rect 30116 29646 30144 31350
rect 30104 29640 30156 29646
rect 30104 29582 30156 29588
rect 29644 29572 29696 29578
rect 29644 29514 29696 29520
rect 29656 29306 29684 29514
rect 29644 29300 29696 29306
rect 29644 29242 29696 29248
rect 29644 29164 29696 29170
rect 29644 29106 29696 29112
rect 29656 28082 29684 29106
rect 29828 29096 29880 29102
rect 29828 29038 29880 29044
rect 29734 28656 29790 28665
rect 29734 28591 29736 28600
rect 29788 28591 29790 28600
rect 29736 28562 29788 28568
rect 29840 28490 29868 29038
rect 29920 28960 29972 28966
rect 29920 28902 29972 28908
rect 29932 28694 29960 28902
rect 29920 28688 29972 28694
rect 29920 28630 29972 28636
rect 30012 28688 30064 28694
rect 30012 28630 30064 28636
rect 29828 28484 29880 28490
rect 29828 28426 29880 28432
rect 29932 28422 29960 28630
rect 30024 28558 30052 28630
rect 30012 28552 30064 28558
rect 30012 28494 30064 28500
rect 29920 28416 29972 28422
rect 29920 28358 29972 28364
rect 29644 28076 29696 28082
rect 29644 28018 29696 28024
rect 29920 28076 29972 28082
rect 29920 28018 29972 28024
rect 29460 27940 29512 27946
rect 29460 27882 29512 27888
rect 29472 27470 29500 27882
rect 29460 27464 29512 27470
rect 29460 27406 29512 27412
rect 29000 27124 29052 27130
rect 29000 27066 29052 27072
rect 29092 27124 29144 27130
rect 29092 27066 29144 27072
rect 28908 27056 28960 27062
rect 29104 27010 29132 27066
rect 28908 26998 28960 27004
rect 29012 26982 29132 27010
rect 29184 26988 29236 26994
rect 29012 26382 29040 26982
rect 29184 26930 29236 26936
rect 29092 26784 29144 26790
rect 29092 26726 29144 26732
rect 29000 26376 29052 26382
rect 29000 26318 29052 26324
rect 29012 25974 29040 26318
rect 29000 25968 29052 25974
rect 29000 25910 29052 25916
rect 28908 25152 28960 25158
rect 28908 25094 28960 25100
rect 28920 24886 28948 25094
rect 28908 24880 28960 24886
rect 28908 24822 28960 24828
rect 29000 24608 29052 24614
rect 29000 24550 29052 24556
rect 28908 24268 28960 24274
rect 28908 24210 28960 24216
rect 28920 22438 28948 24210
rect 29012 23730 29040 24550
rect 29000 23724 29052 23730
rect 29000 23666 29052 23672
rect 28908 22432 28960 22438
rect 28908 22374 28960 22380
rect 28920 22234 28948 22374
rect 28908 22228 28960 22234
rect 28908 22170 28960 22176
rect 28814 22128 28870 22137
rect 28814 22063 28870 22072
rect 28816 22024 28868 22030
rect 28814 21992 28816 22001
rect 28868 21992 28870 22001
rect 28814 21927 28870 21936
rect 28724 20800 28776 20806
rect 28724 20742 28776 20748
rect 28736 20602 28764 20742
rect 28828 20602 28856 21927
rect 29000 21548 29052 21554
rect 29000 21490 29052 21496
rect 29012 20942 29040 21490
rect 29000 20936 29052 20942
rect 29000 20878 29052 20884
rect 28906 20632 28962 20641
rect 28724 20596 28776 20602
rect 28724 20538 28776 20544
rect 28816 20596 28868 20602
rect 28962 20602 29040 20618
rect 28962 20596 29052 20602
rect 28962 20590 29000 20596
rect 28906 20567 28962 20576
rect 28816 20538 28868 20544
rect 29000 20538 29052 20544
rect 28906 20496 28962 20505
rect 28906 20431 28908 20440
rect 28960 20431 28962 20440
rect 28908 20402 28960 20408
rect 29104 20369 29132 26726
rect 29196 25294 29224 26930
rect 29184 25288 29236 25294
rect 29184 25230 29236 25236
rect 29196 24954 29224 25230
rect 29184 24948 29236 24954
rect 29184 24890 29236 24896
rect 29276 22704 29328 22710
rect 29276 22646 29328 22652
rect 29288 21554 29316 22646
rect 29276 21548 29328 21554
rect 29276 21490 29328 21496
rect 29090 20360 29146 20369
rect 28724 20324 28776 20330
rect 28716 20272 28724 20312
rect 29090 20295 29146 20304
rect 28716 20266 28776 20272
rect 28716 20210 28744 20266
rect 29000 20256 29052 20262
rect 28716 20182 28856 20210
rect 29000 20198 29052 20204
rect 29090 20224 29146 20233
rect 28722 20088 28778 20097
rect 28722 20023 28778 20032
rect 28632 17740 28684 17746
rect 28632 17682 28684 17688
rect 28632 17196 28684 17202
rect 28632 17138 28684 17144
rect 28644 16250 28672 17138
rect 28632 16244 28684 16250
rect 28632 16186 28684 16192
rect 28736 16130 28764 20023
rect 28828 19378 28856 20182
rect 29012 20182 29045 20198
rect 29012 19990 29040 20182
rect 29090 20159 29146 20168
rect 29000 19984 29052 19990
rect 29000 19926 29052 19932
rect 28816 19372 28868 19378
rect 28816 19314 28868 19320
rect 28828 17270 28856 19314
rect 28908 17536 28960 17542
rect 28908 17478 28960 17484
rect 28816 17264 28868 17270
rect 28816 17206 28868 17212
rect 28644 16102 28764 16130
rect 28920 16114 28948 17478
rect 28908 16108 28960 16114
rect 28540 16040 28592 16046
rect 28540 15982 28592 15988
rect 28448 15020 28500 15026
rect 28448 14962 28500 14968
rect 28264 14476 28316 14482
rect 28264 14418 28316 14424
rect 28264 14272 28316 14278
rect 28264 14214 28316 14220
rect 28276 13326 28304 14214
rect 28264 13320 28316 13326
rect 28264 13262 28316 13268
rect 28276 12850 28304 13262
rect 28264 12844 28316 12850
rect 28264 12786 28316 12792
rect 28448 12844 28500 12850
rect 28448 12786 28500 12792
rect 28356 12776 28408 12782
rect 28356 12718 28408 12724
rect 28172 12640 28224 12646
rect 28172 12582 28224 12588
rect 28080 7812 28132 7818
rect 28080 7754 28132 7760
rect 27988 7404 28040 7410
rect 27988 7346 28040 7352
rect 27804 7200 27856 7206
rect 27804 7142 27856 7148
rect 28080 6928 28132 6934
rect 28080 6870 28132 6876
rect 28092 6458 28120 6870
rect 28080 6452 28132 6458
rect 28080 6394 28132 6400
rect 27896 5908 27948 5914
rect 27896 5850 27948 5856
rect 27712 5704 27764 5710
rect 27712 5646 27764 5652
rect 27528 5228 27580 5234
rect 27528 5170 27580 5176
rect 27540 4690 27568 5170
rect 27620 5024 27672 5030
rect 27620 4966 27672 4972
rect 27632 4826 27660 4966
rect 27620 4820 27672 4826
rect 27620 4762 27672 4768
rect 27528 4684 27580 4690
rect 27528 4626 27580 4632
rect 27908 4622 27936 5850
rect 27988 5160 28040 5166
rect 27988 5102 28040 5108
rect 28000 4826 28028 5102
rect 27988 4820 28040 4826
rect 27988 4762 28040 4768
rect 27436 4616 27488 4622
rect 27436 4558 27488 4564
rect 27896 4616 27948 4622
rect 27896 4558 27948 4564
rect 27160 4140 27212 4146
rect 27160 4082 27212 4088
rect 27344 4140 27396 4146
rect 27344 4082 27396 4088
rect 27172 3738 27200 4082
rect 27344 4004 27396 4010
rect 27344 3946 27396 3952
rect 27160 3732 27212 3738
rect 27160 3674 27212 3680
rect 27252 3732 27304 3738
rect 27252 3674 27304 3680
rect 27264 800 27292 3674
rect 27356 2378 27384 3946
rect 27344 2372 27396 2378
rect 27344 2314 27396 2320
rect 27448 1426 27476 4558
rect 27528 3936 27580 3942
rect 27528 3878 27580 3884
rect 27620 3936 27672 3942
rect 27620 3878 27672 3884
rect 27540 3777 27568 3878
rect 27526 3768 27582 3777
rect 27526 3703 27582 3712
rect 27436 1420 27488 1426
rect 27436 1362 27488 1368
rect 27632 800 27660 3878
rect 27988 3528 28040 3534
rect 27988 3470 28040 3476
rect 27896 3188 27948 3194
rect 27896 3130 27948 3136
rect 27908 2446 27936 3130
rect 28000 2650 28028 3470
rect 28080 2848 28132 2854
rect 28080 2790 28132 2796
rect 27988 2644 28040 2650
rect 27988 2586 28040 2592
rect 27896 2440 27948 2446
rect 27896 2382 27948 2388
rect 27988 2440 28040 2446
rect 27988 2382 28040 2388
rect 28000 2106 28028 2382
rect 27988 2100 28040 2106
rect 27988 2042 28040 2048
rect 28092 1442 28120 2790
rect 28184 2106 28212 12582
rect 28368 12306 28396 12718
rect 28356 12300 28408 12306
rect 28356 12242 28408 12248
rect 28368 11762 28396 12242
rect 28460 12238 28488 12786
rect 28448 12232 28500 12238
rect 28448 12174 28500 12180
rect 28448 11892 28500 11898
rect 28448 11834 28500 11840
rect 28356 11756 28408 11762
rect 28356 11698 28408 11704
rect 28356 7880 28408 7886
rect 28356 7822 28408 7828
rect 28368 7478 28396 7822
rect 28356 7472 28408 7478
rect 28356 7414 28408 7420
rect 28368 7206 28396 7414
rect 28356 7200 28408 7206
rect 28356 7142 28408 7148
rect 28356 5024 28408 5030
rect 28356 4966 28408 4972
rect 28368 4554 28396 4966
rect 28356 4548 28408 4554
rect 28356 4490 28408 4496
rect 28356 3936 28408 3942
rect 28356 3878 28408 3884
rect 28264 2440 28316 2446
rect 28264 2382 28316 2388
rect 28172 2100 28224 2106
rect 28172 2042 28224 2048
rect 28276 1970 28304 2382
rect 28264 1964 28316 1970
rect 28264 1906 28316 1912
rect 28000 1414 28120 1442
rect 28000 800 28028 1414
rect 28368 800 28396 3878
rect 28460 3641 28488 11834
rect 28644 8090 28672 16102
rect 28908 16050 28960 16056
rect 28816 15496 28868 15502
rect 28816 15438 28868 15444
rect 28724 12640 28776 12646
rect 28724 12582 28776 12588
rect 28736 11898 28764 12582
rect 28828 12238 28856 15438
rect 28920 12850 28948 16050
rect 29000 15020 29052 15026
rect 29000 14962 29052 14968
rect 29012 14618 29040 14962
rect 29000 14612 29052 14618
rect 29000 14554 29052 14560
rect 29104 14482 29132 20159
rect 29288 19334 29316 21490
rect 29368 20392 29420 20398
rect 29368 20334 29420 20340
rect 29380 20262 29408 20334
rect 29368 20256 29420 20262
rect 29368 20198 29420 20204
rect 29472 19334 29500 27406
rect 29552 27328 29604 27334
rect 29552 27270 29604 27276
rect 29564 27062 29592 27270
rect 29552 27056 29604 27062
rect 29552 26998 29604 27004
rect 29552 21616 29604 21622
rect 29550 21584 29552 21593
rect 29604 21584 29606 21593
rect 29550 21519 29606 21528
rect 29656 19334 29684 28018
rect 29932 27606 29960 28018
rect 29920 27600 29972 27606
rect 29920 27542 29972 27548
rect 29736 27532 29788 27538
rect 29736 27474 29788 27480
rect 29748 26314 29776 27474
rect 30012 27464 30064 27470
rect 30012 27406 30064 27412
rect 30024 26586 30052 27406
rect 30116 26790 30144 29582
rect 30288 29164 30340 29170
rect 30288 29106 30340 29112
rect 30300 29034 30328 29106
rect 30196 29028 30248 29034
rect 30196 28970 30248 28976
rect 30288 29028 30340 29034
rect 30288 28970 30340 28976
rect 30208 28558 30236 28970
rect 30196 28552 30248 28558
rect 30196 28494 30248 28500
rect 30392 28150 30420 33594
rect 30484 32026 30512 35158
rect 30576 35086 30604 35702
rect 30840 35692 30892 35698
rect 30840 35634 30892 35640
rect 30748 35488 30800 35494
rect 30748 35430 30800 35436
rect 30564 35080 30616 35086
rect 30564 35022 30616 35028
rect 30760 34202 30788 35430
rect 30852 35018 30880 35634
rect 31036 35290 31064 47126
rect 31496 47054 31524 49286
rect 32034 49286 32352 49314
rect 32034 49200 32090 49286
rect 31484 47048 31536 47054
rect 31484 46990 31536 46996
rect 32324 46578 32352 49286
rect 32862 49200 32918 50000
rect 33690 49314 33746 50000
rect 34518 49314 34574 50000
rect 33690 49286 33916 49314
rect 33690 49200 33746 49286
rect 32404 47048 32456 47054
rect 32404 46990 32456 46996
rect 32312 46572 32364 46578
rect 32312 46514 32364 46520
rect 32128 46368 32180 46374
rect 32128 46310 32180 46316
rect 32140 35562 32168 46310
rect 32128 35556 32180 35562
rect 32128 35498 32180 35504
rect 31024 35284 31076 35290
rect 31024 35226 31076 35232
rect 32416 35154 32444 46990
rect 32876 46578 32904 49200
rect 33888 47054 33916 49286
rect 34518 49286 34744 49314
rect 34518 49200 34574 49286
rect 33876 47048 33928 47054
rect 33876 46990 33928 46996
rect 34060 46980 34112 46986
rect 34060 46922 34112 46928
rect 32864 46572 32916 46578
rect 32864 46514 32916 46520
rect 32956 46368 33008 46374
rect 32956 46310 33008 46316
rect 32968 39642 32996 46310
rect 34072 41274 34100 46922
rect 34716 46646 34744 49286
rect 35346 49200 35402 50000
rect 36174 49314 36230 50000
rect 35912 49286 36230 49314
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 35360 47054 35388 49200
rect 35912 47122 35940 49286
rect 36174 49200 36230 49286
rect 37002 49314 37058 50000
rect 37002 49286 37228 49314
rect 37002 49200 37058 49286
rect 35900 47116 35952 47122
rect 35900 47058 35952 47064
rect 35348 47048 35400 47054
rect 35348 46990 35400 46996
rect 36176 47048 36228 47054
rect 36176 46990 36228 46996
rect 34704 46640 34756 46646
rect 34704 46582 34756 46588
rect 34796 46368 34848 46374
rect 34796 46310 34848 46316
rect 34060 41268 34112 41274
rect 34060 41210 34112 41216
rect 34808 41206 34836 46310
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34796 41200 34848 41206
rect 34796 41142 34848 41148
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 36188 39846 36216 46990
rect 37200 45966 37228 49286
rect 37830 49200 37886 50000
rect 38658 49200 38714 50000
rect 39486 49200 39542 50000
rect 37844 47122 37872 49200
rect 37832 47116 37884 47122
rect 37832 47058 37884 47064
rect 37556 47048 37608 47054
rect 37556 46990 37608 46996
rect 37464 46504 37516 46510
rect 37464 46446 37516 46452
rect 37188 45960 37240 45966
rect 37188 45902 37240 45908
rect 37280 45824 37332 45830
rect 37280 45766 37332 45772
rect 36176 39840 36228 39846
rect 36176 39782 36228 39788
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 32956 39636 33008 39642
rect 32956 39578 33008 39584
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 37292 36378 37320 45766
rect 37476 37738 37504 46446
rect 37464 37732 37516 37738
rect 37464 37674 37516 37680
rect 37280 36372 37332 36378
rect 37280 36314 37332 36320
rect 37568 35630 37596 46990
rect 38672 46578 38700 49200
rect 38660 46572 38712 46578
rect 38660 46514 38712 46520
rect 39500 45966 39528 49200
rect 39488 45960 39540 45966
rect 39488 45902 39540 45908
rect 38016 45824 38068 45830
rect 38016 45766 38068 45772
rect 37556 35624 37608 35630
rect 37556 35566 37608 35572
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 32404 35148 32456 35154
rect 32404 35090 32456 35096
rect 31116 35080 31168 35086
rect 31116 35022 31168 35028
rect 30840 35012 30892 35018
rect 30840 34954 30892 34960
rect 30748 34196 30800 34202
rect 30748 34138 30800 34144
rect 30564 33992 30616 33998
rect 30564 33934 30616 33940
rect 30576 33522 30604 33934
rect 30564 33516 30616 33522
rect 30564 33458 30616 33464
rect 30840 33516 30892 33522
rect 30840 33458 30892 33464
rect 30656 32904 30708 32910
rect 30656 32846 30708 32852
rect 30564 32768 30616 32774
rect 30564 32710 30616 32716
rect 30576 32502 30604 32710
rect 30564 32496 30616 32502
rect 30564 32438 30616 32444
rect 30668 32026 30696 32846
rect 30472 32020 30524 32026
rect 30472 31962 30524 31968
rect 30656 32020 30708 32026
rect 30656 31962 30708 31968
rect 30748 31816 30800 31822
rect 30748 31758 30800 31764
rect 30472 31680 30524 31686
rect 30472 31622 30524 31628
rect 30484 31482 30512 31622
rect 30472 31476 30524 31482
rect 30472 31418 30524 31424
rect 30760 31346 30788 31758
rect 30748 31340 30800 31346
rect 30748 31282 30800 31288
rect 30852 29866 30880 33458
rect 31128 31754 31156 35022
rect 31576 34944 31628 34950
rect 31576 34886 31628 34892
rect 31208 34604 31260 34610
rect 31208 34546 31260 34552
rect 31220 34202 31248 34546
rect 31208 34196 31260 34202
rect 31208 34138 31260 34144
rect 31300 31816 31352 31822
rect 31300 31758 31352 31764
rect 31128 31726 31248 31754
rect 30760 29850 30880 29866
rect 30748 29844 30880 29850
rect 30800 29838 30880 29844
rect 30748 29786 30800 29792
rect 30564 29572 30616 29578
rect 30564 29514 30616 29520
rect 30472 29504 30524 29510
rect 30472 29446 30524 29452
rect 30484 29306 30512 29446
rect 30472 29300 30524 29306
rect 30472 29242 30524 29248
rect 30380 28144 30432 28150
rect 30380 28086 30432 28092
rect 30196 28076 30248 28082
rect 30196 28018 30248 28024
rect 30208 27674 30236 28018
rect 30288 27872 30340 27878
rect 30288 27814 30340 27820
rect 30196 27668 30248 27674
rect 30196 27610 30248 27616
rect 30104 26784 30156 26790
rect 30104 26726 30156 26732
rect 30012 26580 30064 26586
rect 30012 26522 30064 26528
rect 30116 26382 30144 26726
rect 30300 26382 30328 27814
rect 30104 26376 30156 26382
rect 30104 26318 30156 26324
rect 30288 26376 30340 26382
rect 30288 26318 30340 26324
rect 29736 26308 29788 26314
rect 29736 26250 29788 26256
rect 30116 24206 30144 26318
rect 30484 25974 30512 29242
rect 30576 28762 30604 29514
rect 30564 28756 30616 28762
rect 30564 28698 30616 28704
rect 30760 28694 30788 29786
rect 31024 29096 31076 29102
rect 31024 29038 31076 29044
rect 30748 28688 30800 28694
rect 30748 28630 30800 28636
rect 30472 25968 30524 25974
rect 30472 25910 30524 25916
rect 30380 25764 30432 25770
rect 30380 25706 30432 25712
rect 30656 25764 30708 25770
rect 30656 25706 30708 25712
rect 30196 25424 30248 25430
rect 30196 25366 30248 25372
rect 30208 24886 30236 25366
rect 30392 25294 30420 25706
rect 30380 25288 30432 25294
rect 30380 25230 30432 25236
rect 30196 24880 30248 24886
rect 30196 24822 30248 24828
rect 30104 24200 30156 24206
rect 30104 24142 30156 24148
rect 30288 24064 30340 24070
rect 30288 24006 30340 24012
rect 30300 23798 30328 24006
rect 30288 23792 30340 23798
rect 30288 23734 30340 23740
rect 30392 23730 30420 25230
rect 30668 25226 30696 25706
rect 30760 25294 30788 28630
rect 31036 28218 31064 29038
rect 31116 28484 31168 28490
rect 31116 28426 31168 28432
rect 31024 28212 31076 28218
rect 31024 28154 31076 28160
rect 31128 28150 31156 28426
rect 31116 28144 31168 28150
rect 31116 28086 31168 28092
rect 30932 25900 30984 25906
rect 30932 25842 30984 25848
rect 30748 25288 30800 25294
rect 30748 25230 30800 25236
rect 30656 25220 30708 25226
rect 30656 25162 30708 25168
rect 30472 24948 30524 24954
rect 30472 24890 30524 24896
rect 29736 23724 29788 23730
rect 29736 23666 29788 23672
rect 30380 23724 30432 23730
rect 30380 23666 30432 23672
rect 29748 21554 29776 23666
rect 30380 23588 30432 23594
rect 30380 23530 30432 23536
rect 30012 23316 30064 23322
rect 30012 23258 30064 23264
rect 29920 22636 29972 22642
rect 29920 22578 29972 22584
rect 29828 22092 29880 22098
rect 29828 22034 29880 22040
rect 29736 21548 29788 21554
rect 29736 21490 29788 21496
rect 29840 21010 29868 22034
rect 29932 21962 29960 22578
rect 29920 21956 29972 21962
rect 29920 21898 29972 21904
rect 29920 21684 29972 21690
rect 29920 21626 29972 21632
rect 29828 21004 29880 21010
rect 29828 20946 29880 20952
rect 29828 20800 29880 20806
rect 29828 20742 29880 20748
rect 29840 20534 29868 20742
rect 29932 20602 29960 21626
rect 30024 21536 30052 23258
rect 30104 22160 30156 22166
rect 30104 22102 30156 22108
rect 30196 22160 30248 22166
rect 30196 22102 30248 22108
rect 30116 21690 30144 22102
rect 30208 21842 30236 22102
rect 30208 21814 30328 21842
rect 30104 21684 30156 21690
rect 30104 21626 30156 21632
rect 30104 21548 30156 21554
rect 30024 21508 30104 21536
rect 30104 21490 30156 21496
rect 30116 20874 30144 21490
rect 30300 21146 30328 21814
rect 30288 21140 30340 21146
rect 30288 21082 30340 21088
rect 30104 20868 30156 20874
rect 30104 20810 30156 20816
rect 29920 20596 29972 20602
rect 29920 20538 29972 20544
rect 30196 20596 30248 20602
rect 30196 20538 30248 20544
rect 29828 20528 29880 20534
rect 29828 20470 29880 20476
rect 30208 19514 30236 20538
rect 30196 19508 30248 19514
rect 30196 19450 30248 19456
rect 29196 19306 29316 19334
rect 29380 19306 29500 19334
rect 29564 19306 29684 19334
rect 29092 14476 29144 14482
rect 29092 14418 29144 14424
rect 29092 13932 29144 13938
rect 29092 13874 29144 13880
rect 28908 12844 28960 12850
rect 28908 12786 28960 12792
rect 29104 12714 29132 13874
rect 29092 12708 29144 12714
rect 29092 12650 29144 12656
rect 28816 12232 28868 12238
rect 28816 12174 28868 12180
rect 28724 11892 28776 11898
rect 28724 11834 28776 11840
rect 28724 11688 28776 11694
rect 28724 11630 28776 11636
rect 28632 8084 28684 8090
rect 28632 8026 28684 8032
rect 28644 7426 28672 8026
rect 28736 7834 28764 11630
rect 28816 10464 28868 10470
rect 28816 10406 28868 10412
rect 28828 10062 28856 10406
rect 28816 10056 28868 10062
rect 28816 9998 28868 10004
rect 28908 9920 28960 9926
rect 28908 9862 28960 9868
rect 28920 9654 28948 9862
rect 28908 9648 28960 9654
rect 28908 9590 28960 9596
rect 29000 8968 29052 8974
rect 29000 8910 29052 8916
rect 28736 7806 28856 7834
rect 28552 7410 28672 7426
rect 28540 7404 28672 7410
rect 28592 7398 28672 7404
rect 28540 7346 28592 7352
rect 28724 7200 28776 7206
rect 28724 7142 28776 7148
rect 28736 6730 28764 7142
rect 28724 6724 28776 6730
rect 28724 6666 28776 6672
rect 28724 6112 28776 6118
rect 28724 6054 28776 6060
rect 28736 5914 28764 6054
rect 28828 5930 28856 7806
rect 28908 7812 28960 7818
rect 28908 7754 28960 7760
rect 28920 7018 28948 7754
rect 29012 7206 29040 8910
rect 29196 8090 29224 19306
rect 29380 10674 29408 19306
rect 29564 15008 29592 19306
rect 29920 17536 29972 17542
rect 29920 17478 29972 17484
rect 29828 17196 29880 17202
rect 29828 17138 29880 17144
rect 29840 16794 29868 17138
rect 29828 16788 29880 16794
rect 29828 16730 29880 16736
rect 29932 16590 29960 17478
rect 29920 16584 29972 16590
rect 29920 16526 29972 16532
rect 30288 16176 30340 16182
rect 30288 16118 30340 16124
rect 30300 15502 30328 16118
rect 30288 15496 30340 15502
rect 30288 15438 30340 15444
rect 29472 14980 29592 15008
rect 29368 10668 29420 10674
rect 29368 10610 29420 10616
rect 29380 9722 29408 10610
rect 29368 9716 29420 9722
rect 29368 9658 29420 9664
rect 29472 9602 29500 14980
rect 29552 14884 29604 14890
rect 29552 14826 29604 14832
rect 29564 14482 29592 14826
rect 29644 14816 29696 14822
rect 29644 14758 29696 14764
rect 29920 14816 29972 14822
rect 29920 14758 29972 14764
rect 29552 14476 29604 14482
rect 29552 14418 29604 14424
rect 29656 14414 29684 14758
rect 29644 14408 29696 14414
rect 29644 14350 29696 14356
rect 29552 14340 29604 14346
rect 29552 14282 29604 14288
rect 29564 12238 29592 14282
rect 29932 13938 29960 14758
rect 29920 13932 29972 13938
rect 29920 13874 29972 13880
rect 30288 13184 30340 13190
rect 30288 13126 30340 13132
rect 30300 12918 30328 13126
rect 30288 12912 30340 12918
rect 30288 12854 30340 12860
rect 29644 12776 29696 12782
rect 29644 12718 29696 12724
rect 29920 12776 29972 12782
rect 29920 12718 29972 12724
rect 29656 12238 29684 12718
rect 29552 12232 29604 12238
rect 29552 12174 29604 12180
rect 29644 12232 29696 12238
rect 29644 12174 29696 12180
rect 29932 11218 29960 12718
rect 29920 11212 29972 11218
rect 29920 11154 29972 11160
rect 30392 11014 30420 23530
rect 30484 22030 30512 24890
rect 30668 24834 30696 25162
rect 30564 24812 30616 24818
rect 30668 24806 30788 24834
rect 30564 24754 30616 24760
rect 30576 23866 30604 24754
rect 30656 24744 30708 24750
rect 30656 24686 30708 24692
rect 30564 23860 30616 23866
rect 30564 23802 30616 23808
rect 30564 23724 30616 23730
rect 30564 23666 30616 23672
rect 30576 23322 30604 23666
rect 30564 23316 30616 23322
rect 30564 23258 30616 23264
rect 30564 22704 30616 22710
rect 30564 22646 30616 22652
rect 30472 22024 30524 22030
rect 30472 21966 30524 21972
rect 30470 21584 30526 21593
rect 30470 21519 30472 21528
rect 30524 21519 30526 21528
rect 30472 21490 30524 21496
rect 30472 21344 30524 21350
rect 30472 21286 30524 21292
rect 30484 18290 30512 21286
rect 30576 20942 30604 22646
rect 30668 21962 30696 24686
rect 30760 23662 30788 24806
rect 30840 24812 30892 24818
rect 30840 24754 30892 24760
rect 30748 23656 30800 23662
rect 30748 23598 30800 23604
rect 30748 22092 30800 22098
rect 30748 22034 30800 22040
rect 30656 21956 30708 21962
rect 30656 21898 30708 21904
rect 30564 20936 30616 20942
rect 30564 20878 30616 20884
rect 30576 20058 30604 20878
rect 30760 20466 30788 22034
rect 30852 22030 30880 24754
rect 30944 24410 30972 25842
rect 31024 25696 31076 25702
rect 31024 25638 31076 25644
rect 30932 24404 30984 24410
rect 30932 24346 30984 24352
rect 30944 23730 30972 24346
rect 31036 23882 31064 25638
rect 31220 24682 31248 31726
rect 31312 31346 31340 31758
rect 31300 31340 31352 31346
rect 31300 31282 31352 31288
rect 31312 29782 31340 31282
rect 31300 29776 31352 29782
rect 31300 29718 31352 29724
rect 31312 29510 31340 29718
rect 31300 29504 31352 29510
rect 31300 29446 31352 29452
rect 31392 27396 31444 27402
rect 31392 27338 31444 27344
rect 31404 26586 31432 27338
rect 31392 26580 31444 26586
rect 31392 26522 31444 26528
rect 31404 25362 31432 26522
rect 31392 25356 31444 25362
rect 31392 25298 31444 25304
rect 31392 24812 31444 24818
rect 31392 24754 31444 24760
rect 31208 24676 31260 24682
rect 31208 24618 31260 24624
rect 31116 24608 31168 24614
rect 31116 24550 31168 24556
rect 31128 24274 31156 24550
rect 31404 24410 31432 24754
rect 31392 24404 31444 24410
rect 31392 24346 31444 24352
rect 31116 24268 31168 24274
rect 31116 24210 31168 24216
rect 31036 23854 31156 23882
rect 30932 23724 30984 23730
rect 30932 23666 30984 23672
rect 30932 22636 30984 22642
rect 30932 22578 30984 22584
rect 30944 22234 30972 22578
rect 30932 22228 30984 22234
rect 30932 22170 30984 22176
rect 30840 22024 30892 22030
rect 30840 21966 30892 21972
rect 30932 21548 30984 21554
rect 30932 21490 30984 21496
rect 30748 20460 30800 20466
rect 30748 20402 30800 20408
rect 30944 20262 30972 21490
rect 30932 20256 30984 20262
rect 30932 20198 30984 20204
rect 30564 20052 30616 20058
rect 30564 19994 30616 20000
rect 30576 18748 30604 19994
rect 30840 19372 30892 19378
rect 30840 19314 30892 19320
rect 30748 19168 30800 19174
rect 30748 19110 30800 19116
rect 30760 18766 30788 19110
rect 30656 18760 30708 18766
rect 30576 18720 30656 18748
rect 30656 18702 30708 18708
rect 30748 18760 30800 18766
rect 30748 18702 30800 18708
rect 30472 18284 30524 18290
rect 30472 18226 30524 18232
rect 30564 18080 30616 18086
rect 30564 18022 30616 18028
rect 30576 17610 30604 18022
rect 30564 17604 30616 17610
rect 30564 17546 30616 17552
rect 30472 17536 30524 17542
rect 30472 17478 30524 17484
rect 30484 16658 30512 17478
rect 30472 16652 30524 16658
rect 30472 16594 30524 16600
rect 30484 15094 30512 16594
rect 30472 15088 30524 15094
rect 30472 15030 30524 15036
rect 30576 15026 30604 17546
rect 30668 17270 30696 18702
rect 30748 18080 30800 18086
rect 30748 18022 30800 18028
rect 30656 17264 30708 17270
rect 30656 17206 30708 17212
rect 30760 16590 30788 18022
rect 30852 17882 30880 19314
rect 30932 18624 30984 18630
rect 30932 18566 30984 18572
rect 30944 18290 30972 18566
rect 30932 18284 30984 18290
rect 30932 18226 30984 18232
rect 30840 17876 30892 17882
rect 30840 17818 30892 17824
rect 30840 16992 30892 16998
rect 30840 16934 30892 16940
rect 30852 16658 30880 16934
rect 30840 16652 30892 16658
rect 30840 16594 30892 16600
rect 30748 16584 30800 16590
rect 30748 16526 30800 16532
rect 30932 16584 30984 16590
rect 30932 16526 30984 16532
rect 30760 16454 30788 16526
rect 30748 16448 30800 16454
rect 30748 16390 30800 16396
rect 30944 16046 30972 16526
rect 31128 16522 31156 23854
rect 31404 23798 31432 24346
rect 31392 23792 31444 23798
rect 31392 23734 31444 23740
rect 31300 22432 31352 22438
rect 31300 22374 31352 22380
rect 31312 22094 31340 22374
rect 31220 22066 31340 22094
rect 31220 22030 31248 22066
rect 31208 22024 31260 22030
rect 31208 21966 31260 21972
rect 31392 22024 31444 22030
rect 31392 21966 31444 21972
rect 31220 21418 31248 21966
rect 31404 21486 31432 21966
rect 31588 21690 31616 34886
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 31944 29640 31996 29646
rect 31944 29582 31996 29588
rect 31956 28762 31984 29582
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 31944 28756 31996 28762
rect 31944 28698 31996 28704
rect 38028 28665 38056 45766
rect 38014 28656 38070 28665
rect 38014 28591 38070 28600
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 33876 25152 33928 25158
rect 33876 25094 33928 25100
rect 31668 23520 31720 23526
rect 31668 23462 31720 23468
rect 31680 22030 31708 23462
rect 32680 23112 32732 23118
rect 32680 23054 32732 23060
rect 32496 22976 32548 22982
rect 32496 22918 32548 22924
rect 32508 22710 32536 22918
rect 32496 22704 32548 22710
rect 32496 22646 32548 22652
rect 31668 22024 31720 22030
rect 31668 21966 31720 21972
rect 32692 21690 32720 23054
rect 33508 22432 33560 22438
rect 33508 22374 33560 22380
rect 33520 22098 33548 22374
rect 33508 22092 33560 22098
rect 33508 22034 33560 22040
rect 32864 22024 32916 22030
rect 32864 21966 32916 21972
rect 32772 21888 32824 21894
rect 32772 21830 32824 21836
rect 31576 21684 31628 21690
rect 31576 21626 31628 21632
rect 32680 21684 32732 21690
rect 32680 21626 32732 21632
rect 32784 21554 32812 21830
rect 31944 21548 31996 21554
rect 31944 21490 31996 21496
rect 32772 21548 32824 21554
rect 32772 21490 32824 21496
rect 31392 21480 31444 21486
rect 31392 21422 31444 21428
rect 31208 21412 31260 21418
rect 31208 21354 31260 21360
rect 31956 21146 31984 21490
rect 31760 21140 31812 21146
rect 31760 21082 31812 21088
rect 31944 21140 31996 21146
rect 31944 21082 31996 21088
rect 31772 20466 31800 21082
rect 31760 20460 31812 20466
rect 31760 20402 31812 20408
rect 31300 20324 31352 20330
rect 31300 20266 31352 20272
rect 31312 19990 31340 20266
rect 32312 20256 32364 20262
rect 32312 20198 32364 20204
rect 31300 19984 31352 19990
rect 31300 19926 31352 19932
rect 32220 19780 32272 19786
rect 32220 19722 32272 19728
rect 32232 19514 32260 19722
rect 32220 19508 32272 19514
rect 32220 19450 32272 19456
rect 32324 18358 32352 20198
rect 32404 19372 32456 19378
rect 32404 19314 32456 19320
rect 32416 18426 32444 19314
rect 32784 18766 32812 21490
rect 32876 20330 32904 21966
rect 33784 21888 33836 21894
rect 33784 21830 33836 21836
rect 33508 21616 33560 21622
rect 33508 21558 33560 21564
rect 33520 20874 33548 21558
rect 33600 21480 33652 21486
rect 33600 21422 33652 21428
rect 33508 20868 33560 20874
rect 33508 20810 33560 20816
rect 32864 20324 32916 20330
rect 32864 20266 32916 20272
rect 33140 20256 33192 20262
rect 33140 20198 33192 20204
rect 32956 19848 33008 19854
rect 32956 19790 33008 19796
rect 32968 19310 32996 19790
rect 33152 19378 33180 20198
rect 33140 19372 33192 19378
rect 33140 19314 33192 19320
rect 32956 19304 33008 19310
rect 32956 19246 33008 19252
rect 32968 18834 32996 19246
rect 32956 18828 33008 18834
rect 32956 18770 33008 18776
rect 32772 18760 32824 18766
rect 32772 18702 32824 18708
rect 32404 18420 32456 18426
rect 32404 18362 32456 18368
rect 32312 18352 32364 18358
rect 32312 18294 32364 18300
rect 32128 18284 32180 18290
rect 32128 18226 32180 18232
rect 32140 17746 32168 18226
rect 32324 17746 32352 18294
rect 32968 18222 32996 18770
rect 33152 18766 33180 19314
rect 33520 19258 33548 20810
rect 33612 19378 33640 21422
rect 33796 20874 33824 21830
rect 33784 20868 33836 20874
rect 33784 20810 33836 20816
rect 33692 20392 33744 20398
rect 33692 20334 33744 20340
rect 33704 20058 33732 20334
rect 33692 20052 33744 20058
rect 33692 19994 33744 20000
rect 33796 19922 33824 20810
rect 33888 20466 33916 25094
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34152 22636 34204 22642
rect 34152 22578 34204 22584
rect 33968 22432 34020 22438
rect 33968 22374 34020 22380
rect 33980 21622 34008 22374
rect 33968 21616 34020 21622
rect 33968 21558 34020 21564
rect 34164 21146 34192 22578
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34980 22024 35032 22030
rect 34980 21966 35032 21972
rect 34992 21690 35020 21966
rect 34980 21684 35032 21690
rect 34980 21626 35032 21632
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34152 21140 34204 21146
rect 34152 21082 34204 21088
rect 33876 20460 33928 20466
rect 33876 20402 33928 20408
rect 34520 20460 34572 20466
rect 34520 20402 34572 20408
rect 34336 20256 34388 20262
rect 34336 20198 34388 20204
rect 33784 19916 33836 19922
rect 33784 19858 33836 19864
rect 34348 19378 34376 20198
rect 34428 19440 34480 19446
rect 34428 19382 34480 19388
rect 33600 19372 33652 19378
rect 33600 19314 33652 19320
rect 34336 19372 34388 19378
rect 34336 19314 34388 19320
rect 33520 19230 33732 19258
rect 33140 18760 33192 18766
rect 33140 18702 33192 18708
rect 33704 18698 33732 19230
rect 33692 18692 33744 18698
rect 33692 18634 33744 18640
rect 33048 18624 33100 18630
rect 33048 18566 33100 18572
rect 33060 18290 33088 18566
rect 33048 18284 33100 18290
rect 33048 18226 33100 18232
rect 32956 18216 33008 18222
rect 32956 18158 33008 18164
rect 33508 18216 33560 18222
rect 33508 18158 33560 18164
rect 32128 17740 32180 17746
rect 32128 17682 32180 17688
rect 32312 17740 32364 17746
rect 32312 17682 32364 17688
rect 32968 17678 32996 18158
rect 32956 17672 33008 17678
rect 32956 17614 33008 17620
rect 33140 17536 33192 17542
rect 33140 17478 33192 17484
rect 31852 17332 31904 17338
rect 31852 17274 31904 17280
rect 31300 17196 31352 17202
rect 31300 17138 31352 17144
rect 31312 16590 31340 17138
rect 31668 16720 31720 16726
rect 31666 16688 31668 16697
rect 31720 16688 31722 16697
rect 31666 16623 31722 16632
rect 31300 16584 31352 16590
rect 31300 16526 31352 16532
rect 31116 16516 31168 16522
rect 31116 16458 31168 16464
rect 31484 16516 31536 16522
rect 31484 16458 31536 16464
rect 31668 16516 31720 16522
rect 31668 16458 31720 16464
rect 31496 16250 31524 16458
rect 31484 16244 31536 16250
rect 31484 16186 31536 16192
rect 30932 16040 30984 16046
rect 30932 15982 30984 15988
rect 30748 15904 30800 15910
rect 30748 15846 30800 15852
rect 30564 15020 30616 15026
rect 30564 14962 30616 14968
rect 30656 14068 30708 14074
rect 30656 14010 30708 14016
rect 30472 13320 30524 13326
rect 30472 13262 30524 13268
rect 30484 12442 30512 13262
rect 30472 12436 30524 12442
rect 30472 12378 30524 12384
rect 30380 11008 30432 11014
rect 30380 10950 30432 10956
rect 29552 10736 29604 10742
rect 29552 10678 29604 10684
rect 30472 10736 30524 10742
rect 30472 10678 30524 10684
rect 29564 10470 29592 10678
rect 30380 10532 30432 10538
rect 30380 10474 30432 10480
rect 29552 10464 29604 10470
rect 29552 10406 29604 10412
rect 30392 10130 30420 10474
rect 30380 10124 30432 10130
rect 30380 10066 30432 10072
rect 30392 9654 30420 10066
rect 30484 10062 30512 10678
rect 30564 10668 30616 10674
rect 30564 10610 30616 10616
rect 30472 10056 30524 10062
rect 30472 9998 30524 10004
rect 30380 9648 30432 9654
rect 29472 9574 29592 9602
rect 30380 9590 30432 9596
rect 29564 9518 29592 9574
rect 29552 9512 29604 9518
rect 29552 9454 29604 9460
rect 30288 9512 30340 9518
rect 30288 9454 30340 9460
rect 30300 8838 30328 9454
rect 30288 8832 30340 8838
rect 30288 8774 30340 8780
rect 30104 8492 30156 8498
rect 30104 8434 30156 8440
rect 29828 8288 29880 8294
rect 29828 8230 29880 8236
rect 29920 8288 29972 8294
rect 29920 8230 29972 8236
rect 29184 8084 29236 8090
rect 29184 8026 29236 8032
rect 29000 7200 29052 7206
rect 29000 7142 29052 7148
rect 28920 7002 29040 7018
rect 28920 6996 29052 7002
rect 28920 6990 29000 6996
rect 29000 6938 29052 6944
rect 29012 6322 29040 6938
rect 29196 6798 29224 8026
rect 29644 7880 29696 7886
rect 29644 7822 29696 7828
rect 29460 7812 29512 7818
rect 29460 7754 29512 7760
rect 29472 7206 29500 7754
rect 29656 7274 29684 7822
rect 29840 7410 29868 8230
rect 29932 8022 29960 8230
rect 29920 8016 29972 8022
rect 29920 7958 29972 7964
rect 30012 7472 30064 7478
rect 30012 7414 30064 7420
rect 29828 7404 29880 7410
rect 29828 7346 29880 7352
rect 29644 7268 29696 7274
rect 29644 7210 29696 7216
rect 29460 7200 29512 7206
rect 29460 7142 29512 7148
rect 29184 6792 29236 6798
rect 29184 6734 29236 6740
rect 29276 6724 29328 6730
rect 29276 6666 29328 6672
rect 29288 6322 29316 6666
rect 29000 6316 29052 6322
rect 29000 6258 29052 6264
rect 29276 6316 29328 6322
rect 29276 6258 29328 6264
rect 29460 6316 29512 6322
rect 29460 6258 29512 6264
rect 28724 5908 28776 5914
rect 28828 5902 28948 5930
rect 28724 5850 28776 5856
rect 28736 4758 28764 5850
rect 28816 5840 28868 5846
rect 28816 5782 28868 5788
rect 28828 5030 28856 5782
rect 28816 5024 28868 5030
rect 28816 4966 28868 4972
rect 28828 4826 28856 4966
rect 28920 4826 28948 5902
rect 29092 5636 29144 5642
rect 29092 5578 29144 5584
rect 28816 4820 28868 4826
rect 28816 4762 28868 4768
rect 28908 4820 28960 4826
rect 28908 4762 28960 4768
rect 28724 4752 28776 4758
rect 28724 4694 28776 4700
rect 28724 4616 28776 4622
rect 28724 4558 28776 4564
rect 28446 3632 28502 3641
rect 28446 3567 28502 3576
rect 28632 3392 28684 3398
rect 28632 3334 28684 3340
rect 28644 3126 28672 3334
rect 28736 3194 28764 4558
rect 28814 3496 28870 3505
rect 28814 3431 28870 3440
rect 28828 3194 28856 3431
rect 28724 3188 28776 3194
rect 28724 3130 28776 3136
rect 28816 3188 28868 3194
rect 28816 3130 28868 3136
rect 28632 3120 28684 3126
rect 28632 3062 28684 3068
rect 28724 2304 28776 2310
rect 28724 2246 28776 2252
rect 28736 800 28764 2246
rect 29104 800 29132 5578
rect 29472 5137 29500 6258
rect 29552 5568 29604 5574
rect 29552 5510 29604 5516
rect 29458 5128 29514 5137
rect 29458 5063 29514 5072
rect 29460 4480 29512 4486
rect 29460 4422 29512 4428
rect 29472 4078 29500 4422
rect 29564 4282 29592 5510
rect 29656 5302 29684 7210
rect 29920 6792 29972 6798
rect 29920 6734 29972 6740
rect 29932 6322 29960 6734
rect 29920 6316 29972 6322
rect 29920 6258 29972 6264
rect 30024 5914 30052 7414
rect 30116 6662 30144 8434
rect 30288 8424 30340 8430
rect 30288 8366 30340 8372
rect 30300 6798 30328 8366
rect 30380 7404 30432 7410
rect 30380 7346 30432 7352
rect 30288 6792 30340 6798
rect 30288 6734 30340 6740
rect 30104 6656 30156 6662
rect 30104 6598 30156 6604
rect 30392 6458 30420 7346
rect 30472 6656 30524 6662
rect 30472 6598 30524 6604
rect 30380 6452 30432 6458
rect 30380 6394 30432 6400
rect 30484 6322 30512 6598
rect 30472 6316 30524 6322
rect 30472 6258 30524 6264
rect 30012 5908 30064 5914
rect 30012 5850 30064 5856
rect 30576 5846 30604 10610
rect 30564 5840 30616 5846
rect 30564 5782 30616 5788
rect 29920 5704 29972 5710
rect 29920 5646 29972 5652
rect 29736 5568 29788 5574
rect 29736 5510 29788 5516
rect 29644 5296 29696 5302
rect 29644 5238 29696 5244
rect 29656 4622 29684 5238
rect 29644 4616 29696 4622
rect 29644 4558 29696 4564
rect 29552 4276 29604 4282
rect 29552 4218 29604 4224
rect 29460 4072 29512 4078
rect 29460 4014 29512 4020
rect 29552 4072 29604 4078
rect 29552 4014 29604 4020
rect 29564 3346 29592 4014
rect 29472 3318 29592 3346
rect 29472 2378 29500 3318
rect 29656 3058 29684 4558
rect 29644 3052 29696 3058
rect 29644 2994 29696 3000
rect 29748 2774 29776 5510
rect 29828 3936 29880 3942
rect 29828 3878 29880 3884
rect 29840 3670 29868 3878
rect 29932 3738 29960 5646
rect 30380 5568 30432 5574
rect 30380 5510 30432 5516
rect 30392 4214 30420 5510
rect 30472 5228 30524 5234
rect 30472 5170 30524 5176
rect 30380 4208 30432 4214
rect 30380 4150 30432 4156
rect 30378 4040 30434 4049
rect 30378 3975 30380 3984
rect 30432 3975 30434 3984
rect 30380 3946 30432 3952
rect 30484 3942 30512 5170
rect 30564 4480 30616 4486
rect 30564 4422 30616 4428
rect 30472 3936 30524 3942
rect 30472 3878 30524 3884
rect 30576 3754 30604 4422
rect 29920 3732 29972 3738
rect 29920 3674 29972 3680
rect 30288 3732 30340 3738
rect 30288 3674 30340 3680
rect 30392 3726 30604 3754
rect 29828 3664 29880 3670
rect 29828 3606 29880 3612
rect 30012 3528 30064 3534
rect 30012 3470 30064 3476
rect 30196 3528 30248 3534
rect 30196 3470 30248 3476
rect 29828 3460 29880 3466
rect 29828 3402 29880 3408
rect 29564 2746 29776 2774
rect 29460 2372 29512 2378
rect 29460 2314 29512 2320
rect 29564 1442 29592 2746
rect 29472 1414 29592 1442
rect 29472 800 29500 1414
rect 29840 800 29868 3402
rect 30024 3126 30052 3470
rect 30012 3120 30064 3126
rect 30012 3062 30064 3068
rect 30208 2650 30236 3470
rect 30196 2644 30248 2650
rect 30196 2586 30248 2592
rect 30012 2440 30064 2446
rect 30012 2382 30064 2388
rect 30024 1970 30052 2382
rect 30012 1964 30064 1970
rect 30012 1906 30064 1912
rect 30300 1034 30328 3674
rect 30392 2582 30420 3726
rect 30564 3664 30616 3670
rect 30564 3606 30616 3612
rect 30380 2576 30432 2582
rect 30380 2518 30432 2524
rect 30208 1006 30328 1034
rect 30208 800 30236 1006
rect 30576 800 30604 3606
rect 30668 2446 30696 14010
rect 30760 13938 30788 15846
rect 30838 15600 30894 15609
rect 30838 15535 30840 15544
rect 30892 15535 30894 15544
rect 30840 15506 30892 15512
rect 30840 15428 30892 15434
rect 30840 15370 30892 15376
rect 30852 14006 30880 15370
rect 31576 14816 31628 14822
rect 31576 14758 31628 14764
rect 31588 14414 31616 14758
rect 31576 14408 31628 14414
rect 31576 14350 31628 14356
rect 30840 14000 30892 14006
rect 30840 13942 30892 13948
rect 31680 13938 31708 16458
rect 31760 16448 31812 16454
rect 31760 16390 31812 16396
rect 31772 15366 31800 16390
rect 31864 15570 31892 17274
rect 31944 17128 31996 17134
rect 31944 17070 31996 17076
rect 31956 15638 31984 17070
rect 32496 16992 32548 16998
rect 32496 16934 32548 16940
rect 32508 16794 32536 16934
rect 32496 16788 32548 16794
rect 32496 16730 32548 16736
rect 33152 16674 33180 17478
rect 33416 17264 33468 17270
rect 33416 17206 33468 17212
rect 32876 16646 33180 16674
rect 32128 16516 32180 16522
rect 32128 16458 32180 16464
rect 32404 16516 32456 16522
rect 32404 16458 32456 16464
rect 31944 15632 31996 15638
rect 31944 15574 31996 15580
rect 31852 15564 31904 15570
rect 31852 15506 31904 15512
rect 31852 15428 31904 15434
rect 31852 15370 31904 15376
rect 31760 15360 31812 15366
rect 31760 15302 31812 15308
rect 31864 14822 31892 15370
rect 32140 15366 32168 16458
rect 32416 16114 32444 16458
rect 32876 16454 32904 16646
rect 33048 16584 33100 16590
rect 33100 16544 33364 16572
rect 33048 16526 33100 16532
rect 32864 16448 32916 16454
rect 32864 16390 32916 16396
rect 32404 16108 32456 16114
rect 32404 16050 32456 16056
rect 32312 15972 32364 15978
rect 32312 15914 32364 15920
rect 32324 15881 32352 15914
rect 32310 15872 32366 15881
rect 32310 15807 32366 15816
rect 32128 15360 32180 15366
rect 32128 15302 32180 15308
rect 31852 14816 31904 14822
rect 31852 14758 31904 14764
rect 32140 14346 32168 15302
rect 32416 14346 32444 16050
rect 32680 16040 32732 16046
rect 32680 15982 32732 15988
rect 32496 15904 32548 15910
rect 32548 15864 32628 15892
rect 32496 15846 32548 15852
rect 32128 14340 32180 14346
rect 32128 14282 32180 14288
rect 32404 14340 32456 14346
rect 32404 14282 32456 14288
rect 32036 14272 32088 14278
rect 32036 14214 32088 14220
rect 30748 13932 30800 13938
rect 30748 13874 30800 13880
rect 31668 13932 31720 13938
rect 31668 13874 31720 13880
rect 31680 13530 31708 13874
rect 31668 13524 31720 13530
rect 31668 13466 31720 13472
rect 31680 12918 31708 13466
rect 31852 13320 31904 13326
rect 31852 13262 31904 13268
rect 31668 12912 31720 12918
rect 31668 12854 31720 12860
rect 31300 12640 31352 12646
rect 31300 12582 31352 12588
rect 31760 12640 31812 12646
rect 31760 12582 31812 12588
rect 31312 12238 31340 12582
rect 31300 12232 31352 12238
rect 31300 12174 31352 12180
rect 30748 12096 30800 12102
rect 30748 12038 30800 12044
rect 30760 6882 30788 12038
rect 31772 11762 31800 12582
rect 31864 12238 31892 13262
rect 32048 12434 32076 14214
rect 31956 12406 32076 12434
rect 31852 12232 31904 12238
rect 31852 12174 31904 12180
rect 31760 11756 31812 11762
rect 31760 11698 31812 11704
rect 30932 11076 30984 11082
rect 30932 11018 30984 11024
rect 30840 11008 30892 11014
rect 30840 10950 30892 10956
rect 30852 10606 30880 10950
rect 30840 10600 30892 10606
rect 30840 10542 30892 10548
rect 30944 10266 30972 11018
rect 31024 10804 31076 10810
rect 31024 10746 31076 10752
rect 30932 10260 30984 10266
rect 30932 10202 30984 10208
rect 30760 6854 30972 6882
rect 30748 6792 30800 6798
rect 30748 6734 30800 6740
rect 30760 6390 30788 6734
rect 30748 6384 30800 6390
rect 30748 6326 30800 6332
rect 30944 5794 30972 6854
rect 31036 6458 31064 10746
rect 31116 10464 31168 10470
rect 31116 10406 31168 10412
rect 31128 9518 31156 10406
rect 31852 9580 31904 9586
rect 31852 9522 31904 9528
rect 31116 9512 31168 9518
rect 31116 9454 31168 9460
rect 31484 7200 31536 7206
rect 31484 7142 31536 7148
rect 31496 7002 31524 7142
rect 31484 6996 31536 7002
rect 31484 6938 31536 6944
rect 31760 6792 31812 6798
rect 31760 6734 31812 6740
rect 31024 6452 31076 6458
rect 31024 6394 31076 6400
rect 31208 6384 31260 6390
rect 31208 6326 31260 6332
rect 31116 6316 31168 6322
rect 31116 6258 31168 6264
rect 30944 5766 31064 5794
rect 30932 5636 30984 5642
rect 30932 5578 30984 5584
rect 30748 5024 30800 5030
rect 30748 4966 30800 4972
rect 30760 4554 30788 4966
rect 30748 4548 30800 4554
rect 30748 4490 30800 4496
rect 30840 4480 30892 4486
rect 30760 4428 30840 4434
rect 30760 4422 30892 4428
rect 30760 4406 30880 4422
rect 30760 4078 30788 4406
rect 30748 4072 30800 4078
rect 30748 4014 30800 4020
rect 30944 3670 30972 5578
rect 30932 3664 30984 3670
rect 30932 3606 30984 3612
rect 31036 3534 31064 5766
rect 31128 5574 31156 6258
rect 31116 5568 31168 5574
rect 31116 5510 31168 5516
rect 31116 4752 31168 4758
rect 31116 4694 31168 4700
rect 31128 4214 31156 4694
rect 31220 4282 31248 6326
rect 31668 6180 31720 6186
rect 31668 6122 31720 6128
rect 31300 6112 31352 6118
rect 31300 6054 31352 6060
rect 31208 4276 31260 4282
rect 31208 4218 31260 4224
rect 31116 4208 31168 4214
rect 31312 4162 31340 6054
rect 31576 5092 31628 5098
rect 31576 5034 31628 5040
rect 31588 4622 31616 5034
rect 31576 4616 31628 4622
rect 31576 4558 31628 4564
rect 31116 4150 31168 4156
rect 31220 4134 31340 4162
rect 31392 4140 31444 4146
rect 31220 4078 31248 4134
rect 31392 4082 31444 4088
rect 31208 4072 31260 4078
rect 31208 4014 31260 4020
rect 31114 3768 31170 3777
rect 31114 3703 31170 3712
rect 31298 3768 31354 3777
rect 31298 3703 31354 3712
rect 31024 3528 31076 3534
rect 31128 3505 31156 3703
rect 31024 3470 31076 3476
rect 31114 3496 31170 3505
rect 31114 3431 31170 3440
rect 30840 3392 30892 3398
rect 30840 3334 30892 3340
rect 31116 3392 31168 3398
rect 31116 3334 31168 3340
rect 30852 2446 30880 3334
rect 30932 3052 30984 3058
rect 30932 2994 30984 3000
rect 30944 2650 30972 2994
rect 31024 2848 31076 2854
rect 31024 2790 31076 2796
rect 30932 2644 30984 2650
rect 30932 2586 30984 2592
rect 31036 2582 31064 2790
rect 31024 2576 31076 2582
rect 31024 2518 31076 2524
rect 31128 2514 31156 3334
rect 31116 2508 31168 2514
rect 31116 2450 31168 2456
rect 30656 2440 30708 2446
rect 30656 2382 30708 2388
rect 30840 2440 30892 2446
rect 30840 2382 30892 2388
rect 30932 2304 30984 2310
rect 30932 2246 30984 2252
rect 30944 800 30972 2246
rect 31312 800 31340 3703
rect 31404 2922 31432 4082
rect 31484 3936 31536 3942
rect 31484 3878 31536 3884
rect 31392 2916 31444 2922
rect 31392 2858 31444 2864
rect 31496 2378 31524 3878
rect 31588 3058 31616 4558
rect 31680 4214 31708 6122
rect 31668 4208 31720 4214
rect 31668 4150 31720 4156
rect 31668 4072 31720 4078
rect 31668 4014 31720 4020
rect 31680 3777 31708 4014
rect 31666 3768 31722 3777
rect 31666 3703 31722 3712
rect 31772 3448 31800 6734
rect 31864 5234 31892 9522
rect 31956 9466 31984 12406
rect 32140 12170 32168 14282
rect 32600 14006 32628 15864
rect 32692 15502 32720 15982
rect 32680 15496 32732 15502
rect 32680 15438 32732 15444
rect 32692 14958 32720 15438
rect 32864 15360 32916 15366
rect 32864 15302 32916 15308
rect 32876 15162 32904 15302
rect 32864 15156 32916 15162
rect 32864 15098 32916 15104
rect 33140 15156 33192 15162
rect 33140 15098 33192 15104
rect 32680 14952 32732 14958
rect 32680 14894 32732 14900
rect 32680 14476 32732 14482
rect 32680 14418 32732 14424
rect 32588 14000 32640 14006
rect 32588 13942 32640 13948
rect 32692 13938 32720 14418
rect 32772 14340 32824 14346
rect 32772 14282 32824 14288
rect 32680 13932 32732 13938
rect 32680 13874 32732 13880
rect 32784 13190 32812 14282
rect 32864 14068 32916 14074
rect 32864 14010 32916 14016
rect 32876 13258 32904 14010
rect 33152 13938 33180 15098
rect 33336 14634 33364 16544
rect 33428 15162 33456 17206
rect 33416 15156 33468 15162
rect 33416 15098 33468 15104
rect 33336 14606 33456 14634
rect 33428 14278 33456 14606
rect 33324 14272 33376 14278
rect 33324 14214 33376 14220
rect 33416 14272 33468 14278
rect 33416 14214 33468 14220
rect 33140 13932 33192 13938
rect 33140 13874 33192 13880
rect 33336 13326 33364 14214
rect 33324 13320 33376 13326
rect 33324 13262 33376 13268
rect 32864 13252 32916 13258
rect 32864 13194 32916 13200
rect 32772 13184 32824 13190
rect 32772 13126 32824 13132
rect 32588 12436 32640 12442
rect 32588 12378 32640 12384
rect 32128 12164 32180 12170
rect 32128 12106 32180 12112
rect 32600 11694 32628 12378
rect 32784 12306 32812 13126
rect 32772 12300 32824 12306
rect 32772 12242 32824 12248
rect 33232 12164 33284 12170
rect 33232 12106 33284 12112
rect 32588 11688 32640 11694
rect 32588 11630 32640 11636
rect 32600 11286 32628 11630
rect 32588 11280 32640 11286
rect 32588 11222 32640 11228
rect 32404 11144 32456 11150
rect 32404 11086 32456 11092
rect 32036 10056 32088 10062
rect 32036 9998 32088 10004
rect 32048 9654 32076 9998
rect 32036 9648 32088 9654
rect 32036 9590 32088 9596
rect 31956 9438 32076 9466
rect 31944 6248 31996 6254
rect 31944 6190 31996 6196
rect 31956 5302 31984 6190
rect 31944 5296 31996 5302
rect 31944 5238 31996 5244
rect 31852 5228 31904 5234
rect 31852 5170 31904 5176
rect 32048 4978 32076 9438
rect 32220 9376 32272 9382
rect 32220 9318 32272 9324
rect 32232 8906 32260 9318
rect 32220 8900 32272 8906
rect 32220 8842 32272 8848
rect 32312 8492 32364 8498
rect 32312 8434 32364 8440
rect 32324 8022 32352 8434
rect 32312 8016 32364 8022
rect 32312 7958 32364 7964
rect 32416 6882 32444 11086
rect 32600 10606 32628 11222
rect 33244 10810 33272 12106
rect 33324 11552 33376 11558
rect 33324 11494 33376 11500
rect 33232 10804 33284 10810
rect 33232 10746 33284 10752
rect 33336 10742 33364 11494
rect 32772 10736 32824 10742
rect 32772 10678 32824 10684
rect 33324 10736 33376 10742
rect 33324 10678 33376 10684
rect 32588 10600 32640 10606
rect 32588 10542 32640 10548
rect 32600 10062 32628 10542
rect 32680 10192 32732 10198
rect 32680 10134 32732 10140
rect 32588 10056 32640 10062
rect 32588 9998 32640 10004
rect 32600 8974 32628 9998
rect 32588 8968 32640 8974
rect 32588 8910 32640 8916
rect 32600 8430 32628 8910
rect 32588 8424 32640 8430
rect 32588 8366 32640 8372
rect 32600 8022 32628 8366
rect 32588 8016 32640 8022
rect 32588 7958 32640 7964
rect 32692 7954 32720 10134
rect 32680 7948 32732 7954
rect 32680 7890 32732 7896
rect 32680 7200 32732 7206
rect 32680 7142 32732 7148
rect 32324 6866 32444 6882
rect 32312 6860 32444 6866
rect 32364 6854 32444 6860
rect 32312 6802 32364 6808
rect 32128 6792 32180 6798
rect 32128 6734 32180 6740
rect 32140 5574 32168 6734
rect 32324 5710 32352 6802
rect 32692 6798 32720 7142
rect 32680 6792 32732 6798
rect 32680 6734 32732 6740
rect 32784 6458 32812 10678
rect 33140 9172 33192 9178
rect 33140 9114 33192 9120
rect 33152 7750 33180 9114
rect 33232 8288 33284 8294
rect 33232 8230 33284 8236
rect 33244 8090 33272 8230
rect 33232 8084 33284 8090
rect 33232 8026 33284 8032
rect 33140 7744 33192 7750
rect 33140 7686 33192 7692
rect 33152 7478 33180 7686
rect 33140 7472 33192 7478
rect 33140 7414 33192 7420
rect 33244 7426 33272 8026
rect 33520 7562 33548 18158
rect 33704 17610 33732 18634
rect 34440 17678 34468 19382
rect 34532 18970 34560 20402
rect 34796 20392 34848 20398
rect 34796 20334 34848 20340
rect 34808 19514 34836 20334
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 37280 19712 37332 19718
rect 37280 19654 37332 19660
rect 34704 19508 34756 19514
rect 34704 19450 34756 19456
rect 34796 19508 34848 19514
rect 34796 19450 34848 19456
rect 34520 18964 34572 18970
rect 34520 18906 34572 18912
rect 34716 18834 34744 19450
rect 37292 19310 37320 19654
rect 37648 19372 37700 19378
rect 37648 19314 37700 19320
rect 37280 19304 37332 19310
rect 37280 19246 37332 19252
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34704 18828 34756 18834
rect 34704 18770 34756 18776
rect 34980 18760 35032 18766
rect 34980 18702 35032 18708
rect 34520 18216 34572 18222
rect 34992 18193 35020 18702
rect 34520 18158 34572 18164
rect 34978 18184 35034 18193
rect 34532 17882 34560 18158
rect 34978 18119 35034 18128
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34520 17876 34572 17882
rect 34520 17818 34572 17824
rect 34428 17672 34480 17678
rect 34428 17614 34480 17620
rect 33692 17604 33744 17610
rect 33692 17546 33744 17552
rect 34152 17264 34204 17270
rect 34152 17206 34204 17212
rect 33968 17060 34020 17066
rect 33968 17002 34020 17008
rect 33784 16992 33836 16998
rect 33784 16934 33836 16940
rect 33600 16652 33652 16658
rect 33600 16594 33652 16600
rect 33612 13326 33640 16594
rect 33692 16448 33744 16454
rect 33692 16390 33744 16396
rect 33704 15978 33732 16390
rect 33692 15972 33744 15978
rect 33692 15914 33744 15920
rect 33690 15872 33746 15881
rect 33690 15807 33746 15816
rect 33600 13320 33652 13326
rect 33600 13262 33652 13268
rect 33704 13190 33732 15807
rect 33796 15366 33824 16934
rect 33876 15632 33928 15638
rect 33874 15600 33876 15609
rect 33928 15600 33930 15609
rect 33874 15535 33930 15544
rect 33784 15360 33836 15366
rect 33784 15302 33836 15308
rect 33980 14958 34008 17002
rect 33968 14952 34020 14958
rect 33968 14894 34020 14900
rect 34164 13870 34192 17206
rect 34440 17134 34468 17614
rect 36084 17536 36136 17542
rect 36084 17478 36136 17484
rect 34428 17128 34480 17134
rect 34428 17070 34480 17076
rect 34440 16454 34468 17070
rect 34520 16992 34572 16998
rect 34520 16934 34572 16940
rect 34428 16448 34480 16454
rect 34428 16390 34480 16396
rect 34440 16114 34468 16390
rect 34428 16108 34480 16114
rect 34428 16050 34480 16056
rect 34244 15904 34296 15910
rect 34532 15858 34560 16934
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 35808 16788 35860 16794
rect 35808 16730 35860 16736
rect 34796 16652 34848 16658
rect 34796 16594 34848 16600
rect 34704 16516 34756 16522
rect 34704 16458 34756 16464
rect 34612 16108 34664 16114
rect 34612 16050 34664 16056
rect 34296 15852 34560 15858
rect 34244 15846 34560 15852
rect 34256 15830 34560 15846
rect 34428 15496 34480 15502
rect 34428 15438 34480 15444
rect 34244 15428 34296 15434
rect 34244 15370 34296 15376
rect 34256 14074 34284 15370
rect 34440 15026 34468 15438
rect 34520 15360 34572 15366
rect 34520 15302 34572 15308
rect 34428 15020 34480 15026
rect 34428 14962 34480 14968
rect 34440 14482 34468 14962
rect 34428 14476 34480 14482
rect 34428 14418 34480 14424
rect 34244 14068 34296 14074
rect 34244 14010 34296 14016
rect 34440 13938 34468 14418
rect 34532 14346 34560 15302
rect 34624 14618 34652 16050
rect 34612 14612 34664 14618
rect 34612 14554 34664 14560
rect 34520 14340 34572 14346
rect 34520 14282 34572 14288
rect 34428 13932 34480 13938
rect 34428 13874 34480 13880
rect 34612 13932 34664 13938
rect 34612 13874 34664 13880
rect 34152 13864 34204 13870
rect 34152 13806 34204 13812
rect 34624 13530 34652 13874
rect 34716 13734 34744 16458
rect 34808 14414 34836 16594
rect 35716 15904 35768 15910
rect 35716 15846 35768 15852
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34796 14408 34848 14414
rect 34796 14350 34848 14356
rect 35728 14074 35756 15846
rect 35820 15026 35848 16730
rect 35900 15904 35952 15910
rect 35900 15846 35952 15852
rect 35808 15020 35860 15026
rect 35808 14962 35860 14968
rect 35912 14618 35940 15846
rect 35992 15428 36044 15434
rect 35992 15370 36044 15376
rect 35900 14612 35952 14618
rect 35900 14554 35952 14560
rect 35716 14068 35768 14074
rect 35716 14010 35768 14016
rect 34704 13728 34756 13734
rect 34704 13670 34756 13676
rect 34612 13524 34664 13530
rect 34612 13466 34664 13472
rect 34152 13320 34204 13326
rect 34152 13262 34204 13268
rect 33692 13184 33744 13190
rect 33692 13126 33744 13132
rect 34060 12844 34112 12850
rect 34060 12786 34112 12792
rect 33600 12164 33652 12170
rect 33600 12106 33652 12112
rect 33612 10266 33640 12106
rect 33692 12096 33744 12102
rect 33692 12038 33744 12044
rect 33784 12096 33836 12102
rect 33784 12038 33836 12044
rect 33704 11762 33732 12038
rect 33692 11756 33744 11762
rect 33692 11698 33744 11704
rect 33600 10260 33652 10266
rect 33600 10202 33652 10208
rect 33796 10062 33824 12038
rect 34072 11898 34100 12786
rect 34164 12442 34192 13262
rect 34152 12436 34204 12442
rect 34152 12378 34204 12384
rect 34060 11892 34112 11898
rect 34060 11834 34112 11840
rect 34716 11150 34744 13670
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 36004 13530 36032 15370
rect 36096 14414 36124 17478
rect 36450 16688 36506 16697
rect 36450 16623 36506 16632
rect 36464 16114 36492 16623
rect 36544 16448 36596 16454
rect 36544 16390 36596 16396
rect 36452 16108 36504 16114
rect 36452 16050 36504 16056
rect 36556 15570 36584 16390
rect 36544 15564 36596 15570
rect 36544 15506 36596 15512
rect 36084 14408 36136 14414
rect 36084 14350 36136 14356
rect 35992 13524 36044 13530
rect 35992 13466 36044 13472
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 35532 12368 35584 12374
rect 35532 12310 35584 12316
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34704 11144 34756 11150
rect 34704 11086 34756 11092
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 33784 10056 33836 10062
rect 33784 9998 33836 10004
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34612 8900 34664 8906
rect 34612 8842 34664 8848
rect 34624 8498 34652 8842
rect 34612 8492 34664 8498
rect 34612 8434 34664 8440
rect 34796 8492 34848 8498
rect 34796 8434 34848 8440
rect 33968 8356 34020 8362
rect 33968 8298 34020 8304
rect 33980 7886 34008 8298
rect 34520 8288 34572 8294
rect 34520 8230 34572 8236
rect 34532 7886 34560 8230
rect 33968 7880 34020 7886
rect 33968 7822 34020 7828
rect 34520 7880 34572 7886
rect 34520 7822 34572 7828
rect 33520 7534 33640 7562
rect 33244 7398 33456 7426
rect 33140 7336 33192 7342
rect 33140 7278 33192 7284
rect 32772 6452 32824 6458
rect 32772 6394 32824 6400
rect 32956 6316 33008 6322
rect 32956 6258 33008 6264
rect 32404 6248 32456 6254
rect 32404 6190 32456 6196
rect 32312 5704 32364 5710
rect 32312 5646 32364 5652
rect 32128 5568 32180 5574
rect 32128 5510 32180 5516
rect 32140 5166 32168 5510
rect 32128 5160 32180 5166
rect 32128 5102 32180 5108
rect 32416 5030 32444 6190
rect 32968 5930 32996 6258
rect 33152 6118 33180 7278
rect 33324 6656 33376 6662
rect 33324 6598 33376 6604
rect 33336 6322 33364 6598
rect 33324 6316 33376 6322
rect 33324 6258 33376 6264
rect 33428 6186 33456 7398
rect 33416 6180 33468 6186
rect 33416 6122 33468 6128
rect 33140 6112 33192 6118
rect 33140 6054 33192 6060
rect 32968 5902 33180 5930
rect 32404 5024 32456 5030
rect 32048 4950 32168 4978
rect 32404 4966 32456 4972
rect 31852 4480 31904 4486
rect 31852 4422 31904 4428
rect 31864 3534 31892 4422
rect 32036 4276 32088 4282
rect 32036 4218 32088 4224
rect 32048 3534 32076 4218
rect 31852 3528 31904 3534
rect 31852 3470 31904 3476
rect 32036 3528 32088 3534
rect 32036 3470 32088 3476
rect 31680 3420 31800 3448
rect 31576 3052 31628 3058
rect 31576 2994 31628 3000
rect 31484 2372 31536 2378
rect 31484 2314 31536 2320
rect 31680 800 31708 3420
rect 31864 2854 31892 3470
rect 32036 3120 32088 3126
rect 32036 3062 32088 3068
rect 31852 2848 31904 2854
rect 31852 2790 31904 2796
rect 32048 2514 32076 3062
rect 32140 2774 32168 4950
rect 32416 4826 32444 4966
rect 33152 4826 33180 5902
rect 32220 4820 32272 4826
rect 32220 4762 32272 4768
rect 32404 4820 32456 4826
rect 32404 4762 32456 4768
rect 33140 4820 33192 4826
rect 33140 4762 33192 4768
rect 32232 4570 32260 4762
rect 32588 4684 32640 4690
rect 32588 4626 32640 4632
rect 32600 4570 32628 4626
rect 32232 4542 32628 4570
rect 33508 4616 33560 4622
rect 33508 4558 33560 4564
rect 32312 4140 32364 4146
rect 32312 4082 32364 4088
rect 32324 3738 32352 4082
rect 32404 3936 32456 3942
rect 32956 3936 33008 3942
rect 32404 3878 32456 3884
rect 32692 3884 32956 3890
rect 32692 3878 33008 3884
rect 32312 3732 32364 3738
rect 32312 3674 32364 3680
rect 32220 3528 32272 3534
rect 32220 3470 32272 3476
rect 32232 3398 32260 3470
rect 32220 3392 32272 3398
rect 32220 3334 32272 3340
rect 32312 3392 32364 3398
rect 32312 3334 32364 3340
rect 32140 2746 32260 2774
rect 32232 2514 32260 2746
rect 32036 2508 32088 2514
rect 32036 2450 32088 2456
rect 32220 2508 32272 2514
rect 32220 2450 32272 2456
rect 32324 2446 32352 3334
rect 32312 2440 32364 2446
rect 32312 2382 32364 2388
rect 32036 2372 32088 2378
rect 32036 2314 32088 2320
rect 32048 800 32076 2314
rect 32416 800 32444 3878
rect 32692 3862 32996 3878
rect 32692 3602 32720 3862
rect 32772 3732 32824 3738
rect 32772 3674 32824 3680
rect 32680 3596 32732 3602
rect 32680 3538 32732 3544
rect 32784 800 32812 3674
rect 32864 3528 32916 3534
rect 32864 3470 32916 3476
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 32876 3058 32904 3470
rect 32956 3460 33008 3466
rect 32956 3402 33008 3408
rect 32864 3052 32916 3058
rect 32864 2994 32916 3000
rect 32968 2582 32996 3402
rect 33060 2650 33088 3470
rect 33048 2644 33100 2650
rect 33048 2586 33100 2592
rect 32956 2576 33008 2582
rect 32956 2518 33008 2524
rect 33140 2576 33192 2582
rect 33140 2518 33192 2524
rect 33048 2508 33100 2514
rect 33048 2450 33100 2456
rect 33060 2038 33088 2450
rect 33048 2032 33100 2038
rect 33048 1974 33100 1980
rect 33152 800 33180 2518
rect 33520 800 33548 4558
rect 33612 2774 33640 7534
rect 33980 7002 34008 7822
rect 34612 7744 34664 7750
rect 34612 7686 34664 7692
rect 34336 7472 34388 7478
rect 34336 7414 34388 7420
rect 33968 6996 34020 7002
rect 33968 6938 34020 6944
rect 34060 6316 34112 6322
rect 34060 6258 34112 6264
rect 33784 4072 33836 4078
rect 33784 4014 33836 4020
rect 33796 3534 33824 4014
rect 33876 4004 33928 4010
rect 33876 3946 33928 3952
rect 33784 3528 33836 3534
rect 33784 3470 33836 3476
rect 33612 2746 33824 2774
rect 33796 2446 33824 2746
rect 33692 2440 33744 2446
rect 33692 2382 33744 2388
rect 33784 2440 33836 2446
rect 33784 2382 33836 2388
rect 33704 2106 33732 2382
rect 33692 2100 33744 2106
rect 33692 2042 33744 2048
rect 33888 800 33916 3946
rect 34072 3738 34100 6258
rect 34348 4622 34376 7414
rect 34624 7410 34652 7686
rect 34808 7546 34836 8434
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34796 7540 34848 7546
rect 34796 7482 34848 7488
rect 34612 7404 34664 7410
rect 34612 7346 34664 7352
rect 34624 6798 34652 7346
rect 35440 7268 35492 7274
rect 35440 7210 35492 7216
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34612 6792 34664 6798
rect 34612 6734 34664 6740
rect 34796 6656 34848 6662
rect 34796 6598 34848 6604
rect 34704 5908 34756 5914
rect 34704 5850 34756 5856
rect 34520 5636 34572 5642
rect 34520 5578 34572 5584
rect 34532 5370 34560 5578
rect 34520 5364 34572 5370
rect 34520 5306 34572 5312
rect 34612 5228 34664 5234
rect 34612 5170 34664 5176
rect 34336 4616 34388 4622
rect 34336 4558 34388 4564
rect 34348 4282 34376 4558
rect 34428 4548 34480 4554
rect 34428 4490 34480 4496
rect 34336 4276 34388 4282
rect 34336 4218 34388 4224
rect 34060 3732 34112 3738
rect 34060 3674 34112 3680
rect 34348 3466 34376 4218
rect 34440 3534 34468 4490
rect 34520 4480 34572 4486
rect 34520 4422 34572 4428
rect 34532 4146 34560 4422
rect 34624 4282 34652 5170
rect 34716 4622 34744 5850
rect 34704 4616 34756 4622
rect 34704 4558 34756 4564
rect 34612 4276 34664 4282
rect 34612 4218 34664 4224
rect 34520 4140 34572 4146
rect 34520 4082 34572 4088
rect 34612 4140 34664 4146
rect 34612 4082 34664 4088
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 34336 3460 34388 3466
rect 34336 3402 34388 3408
rect 34244 1420 34296 1426
rect 34244 1362 34296 1368
rect 34256 800 34284 1362
rect 34624 800 34652 4082
rect 34808 4049 34836 6598
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 35348 5228 35400 5234
rect 35348 5170 35400 5176
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 35072 4616 35124 4622
rect 35072 4558 35124 4564
rect 35256 4616 35308 4622
rect 35256 4558 35308 4564
rect 35084 4282 35112 4558
rect 35072 4276 35124 4282
rect 35072 4218 35124 4224
rect 34794 4040 34850 4049
rect 35268 4010 35296 4558
rect 34794 3975 34850 3984
rect 35256 4004 35308 4010
rect 35256 3946 35308 3952
rect 34796 3936 34848 3942
rect 34796 3878 34848 3884
rect 34808 3534 34836 3878
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 34704 3528 34756 3534
rect 34704 3470 34756 3476
rect 34796 3528 34848 3534
rect 34796 3470 34848 3476
rect 34716 2854 34744 3470
rect 35164 3460 35216 3466
rect 35164 3402 35216 3408
rect 35176 3194 35204 3402
rect 35256 3392 35308 3398
rect 35256 3334 35308 3340
rect 35164 3188 35216 3194
rect 35164 3130 35216 3136
rect 35268 2990 35296 3334
rect 35256 2984 35308 2990
rect 35256 2926 35308 2932
rect 34704 2848 34756 2854
rect 34704 2790 34756 2796
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 35360 1442 35388 5170
rect 35452 4282 35480 7210
rect 35440 4276 35492 4282
rect 35440 4218 35492 4224
rect 35452 3534 35480 4218
rect 35440 3528 35492 3534
rect 35440 3470 35492 3476
rect 35440 3392 35492 3398
rect 35440 3334 35492 3340
rect 35268 1414 35388 1442
rect 34992 870 35112 898
rect 34992 800 35020 870
rect 23584 734 23796 762
rect 23846 0 23902 800
rect 24214 0 24270 800
rect 24582 0 24638 800
rect 24950 0 25006 800
rect 25318 0 25374 800
rect 25686 0 25742 800
rect 26054 0 26110 800
rect 26422 0 26478 800
rect 26882 0 26938 800
rect 27250 0 27306 800
rect 27618 0 27674 800
rect 27986 0 28042 800
rect 28354 0 28410 800
rect 28722 0 28778 800
rect 29090 0 29146 800
rect 29458 0 29514 800
rect 29826 0 29882 800
rect 30194 0 30250 800
rect 30562 0 30618 800
rect 30930 0 30986 800
rect 31298 0 31354 800
rect 31666 0 31722 800
rect 32034 0 32090 800
rect 32402 0 32458 800
rect 32770 0 32826 800
rect 33138 0 33194 800
rect 33506 0 33562 800
rect 33874 0 33930 800
rect 34242 0 34298 800
rect 34610 0 34666 800
rect 34978 0 35034 800
rect 35084 762 35112 870
rect 35268 762 35296 1414
rect 35452 898 35480 3334
rect 35544 3058 35572 12310
rect 37188 7880 37240 7886
rect 37188 7822 37240 7828
rect 35808 6860 35860 6866
rect 35808 6802 35860 6808
rect 35624 6248 35676 6254
rect 35624 6190 35676 6196
rect 35636 4010 35664 6190
rect 35820 5914 35848 6802
rect 35808 5908 35860 5914
rect 35808 5850 35860 5856
rect 35714 5128 35770 5137
rect 35714 5063 35770 5072
rect 35728 4826 35756 5063
rect 37200 4826 37228 7822
rect 35716 4820 35768 4826
rect 35716 4762 35768 4768
rect 37188 4820 37240 4826
rect 37188 4762 37240 4768
rect 36544 4548 36596 4554
rect 36544 4490 36596 4496
rect 36556 4282 36584 4490
rect 36544 4276 36596 4282
rect 36544 4218 36596 4224
rect 36176 4208 36228 4214
rect 36176 4150 36228 4156
rect 35808 4140 35860 4146
rect 35808 4082 35860 4088
rect 35714 4040 35770 4049
rect 35624 4004 35676 4010
rect 35714 3975 35770 3984
rect 35624 3946 35676 3952
rect 35728 3534 35756 3975
rect 35716 3528 35768 3534
rect 35716 3470 35768 3476
rect 35532 3052 35584 3058
rect 35532 2994 35584 3000
rect 35820 1034 35848 4082
rect 35992 2848 36044 2854
rect 35992 2790 36044 2796
rect 36004 1426 36032 2790
rect 36188 2446 36216 4150
rect 37660 4146 37688 19314
rect 37832 18216 37884 18222
rect 37832 18158 37884 18164
rect 37844 5234 37872 18158
rect 37924 7472 37976 7478
rect 37924 7414 37976 7420
rect 37936 5914 37964 7414
rect 37924 5908 37976 5914
rect 37924 5850 37976 5856
rect 39028 5704 39080 5710
rect 39028 5646 39080 5652
rect 37832 5228 37884 5234
rect 37832 5170 37884 5176
rect 37924 4548 37976 4554
rect 37924 4490 37976 4496
rect 36820 4140 36872 4146
rect 36820 4082 36872 4088
rect 37648 4140 37700 4146
rect 37648 4082 37700 4088
rect 36542 3632 36598 3641
rect 36542 3567 36598 3576
rect 36556 3534 36584 3567
rect 36544 3528 36596 3534
rect 36544 3470 36596 3476
rect 36452 3392 36504 3398
rect 36452 3334 36504 3340
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 36176 2440 36228 2446
rect 36176 2382 36228 2388
rect 35992 1420 36044 1426
rect 35992 1362 36044 1368
rect 35360 870 35480 898
rect 35728 1006 35848 1034
rect 35360 800 35388 870
rect 35728 800 35756 1006
rect 36096 800 36124 2382
rect 36464 800 36492 3334
rect 36832 800 36860 4082
rect 37556 3936 37608 3942
rect 37556 3878 37608 3884
rect 36910 3496 36966 3505
rect 36910 3431 36966 3440
rect 36924 2990 36952 3431
rect 36912 2984 36964 2990
rect 36912 2926 36964 2932
rect 37188 2440 37240 2446
rect 37188 2382 37240 2388
rect 37200 800 37228 2382
rect 37568 800 37596 3878
rect 37936 800 37964 4490
rect 38660 4480 38712 4486
rect 38660 4422 38712 4428
rect 38292 3052 38344 3058
rect 38292 2994 38344 3000
rect 38304 800 38332 2994
rect 38672 800 38700 4422
rect 39040 800 39068 5646
rect 39764 5024 39816 5030
rect 39764 4966 39816 4972
rect 39396 3460 39448 3466
rect 39396 3402 39448 3408
rect 39408 800 39436 3402
rect 39776 800 39804 4966
rect 35084 734 35296 762
rect 35346 0 35402 800
rect 35714 0 35770 800
rect 36082 0 36138 800
rect 36450 0 36506 800
rect 36818 0 36874 800
rect 37186 0 37242 800
rect 37554 0 37610 800
rect 37922 0 37978 800
rect 38290 0 38346 800
rect 38658 0 38714 800
rect 39026 0 39082 800
rect 39394 0 39450 800
rect 39762 0 39818 800
<< via2 >>
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 10322 37068 10324 37088
rect 10324 37068 10376 37088
rect 10376 37068 10378 37088
rect 10322 37032 10378 37068
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 11150 35128 11206 35184
rect 12530 35672 12586 35728
rect 12346 33224 12402 33280
rect 12346 29180 12348 29200
rect 12348 29180 12400 29200
rect 12400 29180 12402 29200
rect 12346 29144 12402 29180
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 5262 15816 5318 15872
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 1950 2508 2006 2544
rect 1950 2488 1952 2508
rect 1952 2488 2004 2508
rect 2004 2488 2006 2508
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 7286 15852 7288 15872
rect 7288 15852 7340 15872
rect 7340 15852 7342 15872
rect 7286 15816 7342 15852
rect 9402 17448 9458 17504
rect 8206 8084 8262 8120
rect 8206 8064 8208 8084
rect 8208 8064 8260 8084
rect 8260 8064 8262 8084
rect 11334 16652 11390 16688
rect 11334 16632 11336 16652
rect 11336 16632 11388 16652
rect 11388 16632 11390 16652
rect 9632 3596 9688 3598
rect 9632 3544 9634 3596
rect 9634 3544 9686 3596
rect 9686 3544 9688 3596
rect 9632 3542 9688 3544
rect 9770 3460 9826 3496
rect 9770 3440 9772 3460
rect 9772 3440 9824 3460
rect 9824 3440 9826 3460
rect 10690 3440 10746 3496
rect 11150 6724 11206 6760
rect 11150 6704 11152 6724
rect 11152 6704 11204 6724
rect 11204 6704 11206 6724
rect 11518 3576 11574 3632
rect 12990 35128 13046 35184
rect 12714 29144 12770 29200
rect 13450 41248 13506 41304
rect 13726 40704 13782 40760
rect 13174 27104 13230 27160
rect 13634 33516 13690 33552
rect 13634 33496 13636 33516
rect 13636 33496 13688 33516
rect 13688 33496 13690 33516
rect 13358 25780 13360 25800
rect 13360 25780 13412 25800
rect 13412 25780 13414 25800
rect 13358 25744 13414 25780
rect 12898 17992 12954 18048
rect 12806 12688 12862 12744
rect 12898 6724 12954 6760
rect 12898 6704 12900 6724
rect 12900 6704 12952 6724
rect 12952 6704 12954 6724
rect 14278 33260 14280 33280
rect 14280 33260 14332 33280
rect 14332 33260 14334 33280
rect 14278 33224 14334 33260
rect 14186 28908 14188 28928
rect 14188 28908 14240 28928
rect 14240 28908 14242 28928
rect 14186 28872 14242 28908
rect 13910 23568 13966 23624
rect 14278 23568 14334 23624
rect 14922 33516 14978 33552
rect 14922 33496 14924 33516
rect 14924 33496 14976 33516
rect 14976 33496 14978 33516
rect 15566 40976 15622 41032
rect 15382 40840 15438 40896
rect 15842 41148 15844 41168
rect 15844 41148 15896 41168
rect 15896 41148 15898 41168
rect 15842 41112 15898 41148
rect 15934 40976 15990 41032
rect 14922 33224 14978 33280
rect 14278 12688 14334 12744
rect 16486 40840 16542 40896
rect 16394 40704 16450 40760
rect 14922 21548 14978 21584
rect 14922 21528 14924 21548
rect 14924 21528 14976 21548
rect 14976 21528 14978 21548
rect 14922 20460 14978 20496
rect 14922 20440 14924 20460
rect 14924 20440 14976 20460
rect 14976 20440 14978 20460
rect 15290 20304 15346 20360
rect 16026 37324 16082 37360
rect 16026 37304 16028 37324
rect 16028 37304 16080 37324
rect 16080 37304 16082 37324
rect 16026 28872 16082 28928
rect 15566 20304 15622 20360
rect 15290 16632 15346 16688
rect 16486 21564 16488 21584
rect 16488 21564 16540 21584
rect 16540 21564 16542 21584
rect 16486 21528 16542 21564
rect 17682 37324 17738 37360
rect 17682 37304 17684 37324
rect 17684 37304 17736 37324
rect 17736 37304 17738 37324
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 18326 41268 18382 41304
rect 18326 41248 18328 41268
rect 18328 41248 18380 41268
rect 18380 41248 18382 41268
rect 18234 41148 18236 41168
rect 18236 41148 18288 41168
rect 18288 41148 18290 41168
rect 18234 41112 18290 41148
rect 18326 40976 18382 41032
rect 17774 37032 17830 37088
rect 17130 35672 17186 35728
rect 17222 27124 17278 27160
rect 17222 27104 17224 27124
rect 17224 27104 17276 27124
rect 17276 27104 17278 27124
rect 16210 16632 16266 16688
rect 14554 12280 14610 12336
rect 15014 12280 15070 12336
rect 14646 4256 14702 4312
rect 16486 14492 16488 14512
rect 16488 14492 16540 14512
rect 16540 14492 16542 14512
rect 16486 14456 16542 14492
rect 15198 3984 15254 4040
rect 17590 18128 17646 18184
rect 17590 16532 17592 16552
rect 17592 16532 17644 16552
rect 17644 16532 17646 16552
rect 17590 16496 17646 16532
rect 17958 32000 18014 32056
rect 18234 32000 18290 32056
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 17038 4256 17094 4312
rect 18326 18536 18382 18592
rect 18326 14456 18382 14512
rect 19062 34040 19118 34096
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 20074 34448 20130 34504
rect 20074 34060 20130 34096
rect 20074 34040 20076 34060
rect 20076 34040 20128 34060
rect 20128 34040 20130 34060
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19706 32852 19708 32872
rect 19708 32852 19760 32872
rect 19760 32852 19762 32872
rect 19706 32816 19762 32852
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19430 29824 19486 29880
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19798 28620 19854 28656
rect 19798 28600 19800 28620
rect 19800 28600 19852 28620
rect 19852 28600 19854 28620
rect 19706 28500 19708 28520
rect 19708 28500 19760 28520
rect 19760 28500 19762 28520
rect 19706 28464 19762 28500
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19338 27648 19394 27704
rect 19338 27376 19394 27432
rect 19890 28056 19946 28112
rect 19522 27920 19578 27976
rect 19890 27376 19946 27432
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 18602 18148 18658 18184
rect 18602 18128 18604 18148
rect 18604 18128 18656 18148
rect 18656 18128 18658 18148
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19706 25356 19762 25392
rect 19706 25336 19708 25356
rect 19708 25336 19760 25356
rect 19760 25336 19762 25356
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19522 24248 19578 24304
rect 19338 24112 19394 24168
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19338 23704 19394 23760
rect 19522 23740 19524 23760
rect 19524 23740 19576 23760
rect 19576 23740 19578 23760
rect 19522 23704 19578 23740
rect 19154 23568 19210 23624
rect 20442 34584 20498 34640
rect 20350 34484 20352 34504
rect 20352 34484 20404 34504
rect 20404 34484 20406 34504
rect 20350 34448 20406 34484
rect 20534 34040 20590 34096
rect 20442 32816 20498 32872
rect 20442 28464 20498 28520
rect 20534 28328 20590 28384
rect 19062 18808 19118 18864
rect 18878 18672 18934 18728
rect 18970 18400 19026 18456
rect 18878 12280 18934 12336
rect 18602 6840 18658 6896
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 20074 20460 20130 20496
rect 20074 20440 20076 20460
rect 20076 20440 20128 20460
rect 20128 20440 20130 20460
rect 20258 23160 20314 23216
rect 19982 18944 20038 19000
rect 19522 18672 19578 18728
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 20074 18536 20130 18592
rect 19982 17992 20038 18048
rect 19890 17856 19946 17912
rect 19706 17720 19762 17776
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19522 17196 19578 17232
rect 19522 17176 19524 17196
rect 19524 17176 19576 17196
rect 19576 17176 19578 17196
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19706 15428 19762 15464
rect 19706 15408 19708 15428
rect 19708 15408 19760 15428
rect 19760 15408 19762 15428
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 20166 17196 20222 17232
rect 20166 17176 20168 17196
rect 20168 17176 20220 17196
rect 20220 17176 20222 17196
rect 20074 17040 20130 17096
rect 20166 15136 20222 15192
rect 19798 12436 19854 12472
rect 19798 12416 19800 12436
rect 19800 12416 19852 12436
rect 19852 12416 19854 12436
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 20166 12144 20222 12200
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 20442 24248 20498 24304
rect 20994 37204 20996 37224
rect 20996 37204 21048 37224
rect 21048 37204 21050 37224
rect 20994 37168 21050 37204
rect 20718 27512 20774 27568
rect 20902 27920 20958 27976
rect 20626 24132 20682 24168
rect 20626 24112 20628 24132
rect 20628 24112 20680 24132
rect 20680 24112 20682 24132
rect 20442 20032 20498 20088
rect 20350 17992 20406 18048
rect 22006 41132 22062 41168
rect 22006 41112 22008 41132
rect 22008 41112 22060 41132
rect 22060 41112 22062 41132
rect 22282 41148 22284 41168
rect 22284 41148 22336 41168
rect 22336 41148 22338 41168
rect 22282 41112 22338 41148
rect 22006 38412 22062 38448
rect 22006 38392 22008 38412
rect 22008 38392 22060 38412
rect 22060 38392 22062 38412
rect 21362 27512 21418 27568
rect 21178 25336 21234 25392
rect 20810 18400 20866 18456
rect 20718 18128 20774 18184
rect 20718 17992 20774 18048
rect 20810 17856 20866 17912
rect 20718 17176 20774 17232
rect 20442 15408 20498 15464
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19522 6740 19524 6760
rect 19524 6740 19576 6760
rect 19576 6740 19578 6760
rect 19522 6704 19578 6740
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19706 4664 19762 4720
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19890 3440 19946 3496
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20626 12144 20682 12200
rect 21086 18264 21142 18320
rect 21086 6704 21142 6760
rect 20810 4800 20866 4856
rect 21362 20440 21418 20496
rect 21270 18264 21326 18320
rect 21822 28464 21878 28520
rect 22006 28464 22062 28520
rect 22006 23840 22062 23896
rect 22742 32852 22744 32872
rect 22744 32852 22796 32872
rect 22796 32852 22798 32872
rect 22742 32816 22798 32852
rect 22650 28600 22706 28656
rect 22926 28056 22982 28112
rect 23294 29588 23296 29608
rect 23296 29588 23348 29608
rect 23348 29588 23350 29608
rect 23294 29552 23350 29588
rect 23570 27376 23626 27432
rect 22742 21800 22798 21856
rect 21270 8472 21326 8528
rect 22190 8472 22246 8528
rect 21730 4684 21786 4720
rect 21730 4664 21732 4684
rect 21732 4664 21784 4684
rect 21784 4664 21786 4684
rect 22006 4820 22062 4856
rect 22006 4800 22008 4820
rect 22008 4800 22060 4820
rect 22060 4800 22062 4820
rect 23754 28872 23810 28928
rect 24490 34040 24546 34096
rect 23662 21936 23718 21992
rect 24306 27648 24362 27704
rect 25318 38392 25374 38448
rect 24950 29552 25006 29608
rect 24674 23840 24730 23896
rect 23294 17040 23350 17096
rect 25134 29008 25190 29064
rect 25778 32816 25834 32872
rect 26422 37168 26478 37224
rect 25134 21800 25190 21856
rect 24766 19624 24822 19680
rect 24674 17720 24730 17776
rect 23938 4684 23994 4720
rect 23938 4664 23940 4684
rect 23940 4664 23992 4684
rect 23992 4664 23994 4684
rect 28078 29008 28134 29064
rect 25686 24112 25742 24168
rect 25410 20460 25466 20496
rect 25410 20440 25412 20460
rect 25412 20440 25464 20460
rect 25464 20440 25466 20460
rect 25686 20848 25742 20904
rect 24950 6840 25006 6896
rect 26146 21800 26202 21856
rect 26238 9560 26294 9616
rect 27434 20440 27490 20496
rect 27342 19760 27398 19816
rect 27802 27240 27858 27296
rect 27710 25236 27712 25256
rect 27712 25236 27764 25256
rect 27764 25236 27766 25256
rect 27710 25200 27766 25236
rect 27710 21684 27766 21720
rect 27710 21664 27712 21684
rect 27712 21664 27764 21684
rect 27764 21664 27766 21684
rect 27710 21528 27766 21584
rect 27894 21664 27950 21720
rect 27894 21548 27950 21584
rect 27894 21528 27896 21548
rect 27896 21528 27948 21548
rect 27948 21528 27950 21548
rect 28262 27412 28264 27432
rect 28264 27412 28316 27432
rect 28316 27412 28318 27432
rect 28262 27376 28318 27412
rect 28354 27240 28410 27296
rect 28078 22480 28134 22536
rect 28354 22480 28410 22536
rect 28078 20868 28134 20904
rect 28078 20848 28080 20868
rect 28080 20848 28132 20868
rect 28132 20848 28134 20868
rect 28078 20576 28134 20632
rect 27526 9560 27582 9616
rect 28446 20440 28502 20496
rect 28354 19780 28410 19816
rect 28354 19760 28356 19780
rect 28356 19760 28408 19780
rect 28408 19760 28410 19780
rect 28446 19624 28502 19680
rect 29734 28620 29790 28656
rect 29734 28600 29736 28620
rect 29736 28600 29788 28620
rect 29788 28600 29790 28620
rect 28814 22072 28870 22128
rect 28814 21972 28816 21992
rect 28816 21972 28868 21992
rect 28868 21972 28870 21992
rect 28814 21936 28870 21972
rect 28906 20576 28962 20632
rect 28906 20460 28962 20496
rect 28906 20440 28908 20460
rect 28908 20440 28960 20460
rect 28960 20440 28962 20460
rect 29090 20304 29146 20360
rect 28722 20032 28778 20088
rect 29090 20168 29146 20224
rect 27526 3712 27582 3768
rect 29550 21564 29552 21584
rect 29552 21564 29604 21584
rect 29604 21564 29606 21584
rect 29550 21528 29606 21564
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 30470 21548 30526 21584
rect 30470 21528 30472 21548
rect 30472 21528 30524 21548
rect 30524 21528 30526 21548
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 38014 28600 38070 28656
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 31666 16668 31668 16688
rect 31668 16668 31720 16688
rect 31720 16668 31722 16688
rect 31666 16632 31722 16668
rect 28446 3576 28502 3632
rect 28814 3440 28870 3496
rect 29458 5072 29514 5128
rect 30378 4004 30434 4040
rect 30378 3984 30380 4004
rect 30380 3984 30432 4004
rect 30432 3984 30434 4004
rect 30838 15564 30894 15600
rect 30838 15544 30840 15564
rect 30840 15544 30892 15564
rect 30892 15544 30894 15564
rect 32310 15816 32366 15872
rect 31114 3712 31170 3768
rect 31298 3712 31354 3768
rect 31114 3440 31170 3496
rect 31666 3712 31722 3768
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34978 18128 35034 18184
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 33690 15816 33746 15872
rect 33874 15580 33876 15600
rect 33876 15580 33928 15600
rect 33928 15580 33930 15600
rect 33874 15544 33930 15580
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 36450 16632 36506 16688
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34794 3984 34850 4040
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35714 5072 35770 5128
rect 35714 3984 35770 4040
rect 36542 3576 36598 3632
rect 36910 3440 36966 3496
<< metal3 >>
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 13445 41306 13511 41309
rect 18321 41306 18387 41309
rect 13445 41304 18387 41306
rect 13445 41248 13450 41304
rect 13506 41248 18326 41304
rect 18382 41248 18387 41304
rect 13445 41246 18387 41248
rect 13445 41243 13511 41246
rect 18321 41243 18387 41246
rect 15837 41170 15903 41173
rect 18229 41170 18295 41173
rect 15837 41168 18295 41170
rect 15837 41112 15842 41168
rect 15898 41112 18234 41168
rect 18290 41112 18295 41168
rect 15837 41110 18295 41112
rect 15837 41107 15903 41110
rect 18229 41107 18295 41110
rect 22001 41170 22067 41173
rect 22277 41170 22343 41173
rect 22001 41168 22343 41170
rect 22001 41112 22006 41168
rect 22062 41112 22282 41168
rect 22338 41112 22343 41168
rect 22001 41110 22343 41112
rect 22001 41107 22067 41110
rect 22277 41107 22343 41110
rect 15561 41034 15627 41037
rect 15929 41034 15995 41037
rect 18321 41034 18387 41037
rect 15561 41032 18387 41034
rect 15561 40976 15566 41032
rect 15622 40976 15934 41032
rect 15990 40976 18326 41032
rect 18382 40976 18387 41032
rect 15561 40974 18387 40976
rect 15561 40971 15627 40974
rect 15929 40971 15995 40974
rect 18321 40971 18387 40974
rect 15377 40898 15443 40901
rect 16481 40898 16547 40901
rect 15377 40896 16547 40898
rect 15377 40840 15382 40896
rect 15438 40840 16486 40896
rect 16542 40840 16547 40896
rect 15377 40838 16547 40840
rect 15377 40835 15443 40838
rect 16481 40835 16547 40838
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 13721 40762 13787 40765
rect 16389 40762 16455 40765
rect 13721 40760 16455 40762
rect 13721 40704 13726 40760
rect 13782 40704 16394 40760
rect 16450 40704 16455 40760
rect 13721 40702 16455 40704
rect 13721 40699 13787 40702
rect 16389 40699 16455 40702
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 22001 38450 22067 38453
rect 25313 38450 25379 38453
rect 22001 38448 25379 38450
rect 22001 38392 22006 38448
rect 22062 38392 25318 38448
rect 25374 38392 25379 38448
rect 22001 38390 25379 38392
rect 22001 38387 22067 38390
rect 25313 38387 25379 38390
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 16021 37364 16087 37365
rect 17677 37364 17743 37365
rect 16021 37360 16068 37364
rect 16132 37362 16138 37364
rect 16021 37304 16026 37360
rect 16021 37300 16068 37304
rect 16132 37302 16178 37362
rect 17677 37360 17724 37364
rect 17788 37362 17794 37364
rect 17677 37304 17682 37360
rect 16132 37300 16138 37302
rect 17677 37300 17724 37304
rect 17788 37302 17834 37362
rect 17788 37300 17794 37302
rect 16021 37299 16087 37300
rect 17677 37299 17743 37300
rect 20989 37226 21055 37229
rect 26417 37226 26483 37229
rect 20989 37224 26483 37226
rect 20989 37168 20994 37224
rect 21050 37168 26422 37224
rect 26478 37168 26483 37224
rect 20989 37166 26483 37168
rect 20989 37163 21055 37166
rect 26417 37163 26483 37166
rect 10317 37090 10383 37093
rect 17769 37090 17835 37093
rect 10317 37088 17835 37090
rect 10317 37032 10322 37088
rect 10378 37032 17774 37088
rect 17830 37032 17835 37088
rect 10317 37030 17835 37032
rect 10317 37027 10383 37030
rect 17769 37027 17835 37030
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 12525 35730 12591 35733
rect 17125 35730 17191 35733
rect 12525 35728 17191 35730
rect 12525 35672 12530 35728
rect 12586 35672 17130 35728
rect 17186 35672 17191 35728
rect 12525 35670 17191 35672
rect 12525 35667 12591 35670
rect 17125 35667 17191 35670
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 11145 35186 11211 35189
rect 12985 35186 13051 35189
rect 11145 35184 13051 35186
rect 11145 35128 11150 35184
rect 11206 35128 12990 35184
rect 13046 35128 13051 35184
rect 11145 35126 13051 35128
rect 11145 35123 11211 35126
rect 12985 35123 13051 35126
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 20110 34580 20116 34644
rect 20180 34642 20186 34644
rect 20437 34642 20503 34645
rect 20180 34640 20503 34642
rect 20180 34584 20442 34640
rect 20498 34584 20503 34640
rect 20180 34582 20503 34584
rect 20180 34580 20186 34582
rect 20437 34579 20503 34582
rect 20069 34506 20135 34509
rect 20345 34506 20411 34509
rect 20069 34504 20411 34506
rect 20069 34448 20074 34504
rect 20130 34448 20350 34504
rect 20406 34448 20411 34504
rect 20069 34446 20411 34448
rect 20069 34443 20135 34446
rect 20345 34443 20411 34446
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 19057 34098 19123 34101
rect 20069 34098 20135 34101
rect 19057 34096 20135 34098
rect 19057 34040 19062 34096
rect 19118 34040 20074 34096
rect 20130 34040 20135 34096
rect 19057 34038 20135 34040
rect 19057 34035 19123 34038
rect 20069 34035 20135 34038
rect 20529 34098 20595 34101
rect 24485 34098 24551 34101
rect 20529 34096 24551 34098
rect 20529 34040 20534 34096
rect 20590 34040 24490 34096
rect 24546 34040 24551 34096
rect 20529 34038 24551 34040
rect 20529 34035 20595 34038
rect 24485 34035 24551 34038
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 13629 33554 13695 33557
rect 14917 33554 14983 33557
rect 13629 33552 14983 33554
rect 13629 33496 13634 33552
rect 13690 33496 14922 33552
rect 14978 33496 14983 33552
rect 13629 33494 14983 33496
rect 13629 33491 13695 33494
rect 14917 33491 14983 33494
rect 12341 33282 12407 33285
rect 14273 33282 14339 33285
rect 14917 33282 14983 33285
rect 12341 33280 14983 33282
rect 12341 33224 12346 33280
rect 12402 33224 14278 33280
rect 14334 33224 14922 33280
rect 14978 33224 14983 33280
rect 12341 33222 14983 33224
rect 12341 33219 12407 33222
rect 14273 33219 14339 33222
rect 14917 33219 14983 33222
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 19701 32874 19767 32877
rect 20437 32874 20503 32877
rect 22737 32874 22803 32877
rect 25773 32874 25839 32877
rect 19701 32872 25839 32874
rect 19701 32816 19706 32872
rect 19762 32816 20442 32872
rect 20498 32816 22742 32872
rect 22798 32816 25778 32872
rect 25834 32816 25839 32872
rect 19701 32814 25839 32816
rect 19701 32811 19767 32814
rect 20437 32811 20503 32814
rect 22737 32811 22803 32814
rect 25773 32811 25839 32814
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 17953 32058 18019 32061
rect 18229 32058 18295 32061
rect 17953 32056 18295 32058
rect 17953 32000 17958 32056
rect 18014 32000 18234 32056
rect 18290 32000 18295 32056
rect 17953 31998 18295 32000
rect 17953 31995 18019 31998
rect 18229 31995 18295 31998
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 19425 29882 19491 29885
rect 20110 29882 20116 29884
rect 19425 29880 20116 29882
rect 19425 29824 19430 29880
rect 19486 29824 20116 29880
rect 19425 29822 20116 29824
rect 19425 29819 19491 29822
rect 20110 29820 20116 29822
rect 20180 29820 20186 29884
rect 23289 29610 23355 29613
rect 24945 29610 25011 29613
rect 23289 29608 25011 29610
rect 23289 29552 23294 29608
rect 23350 29552 24950 29608
rect 25006 29552 25011 29608
rect 23289 29550 25011 29552
rect 23289 29547 23355 29550
rect 24945 29547 25011 29550
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 12341 29202 12407 29205
rect 12709 29202 12775 29205
rect 12341 29200 12775 29202
rect 12341 29144 12346 29200
rect 12402 29144 12714 29200
rect 12770 29144 12775 29200
rect 12341 29142 12775 29144
rect 12341 29139 12407 29142
rect 12709 29139 12775 29142
rect 25129 29066 25195 29069
rect 28073 29066 28139 29069
rect 25129 29064 28139 29066
rect 25129 29008 25134 29064
rect 25190 29008 28078 29064
rect 28134 29008 28139 29064
rect 25129 29006 28139 29008
rect 25129 29003 25195 29006
rect 28073 29003 28139 29006
rect 14181 28930 14247 28933
rect 16021 28930 16087 28933
rect 23749 28930 23815 28933
rect 14181 28928 23815 28930
rect 14181 28872 14186 28928
rect 14242 28872 16026 28928
rect 16082 28872 23754 28928
rect 23810 28872 23815 28928
rect 14181 28870 23815 28872
rect 14181 28867 14247 28870
rect 16021 28867 16087 28870
rect 23749 28867 23815 28870
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 19793 28658 19859 28661
rect 20294 28658 20300 28660
rect 19793 28656 20300 28658
rect 19793 28600 19798 28656
rect 19854 28600 20300 28656
rect 19793 28598 20300 28600
rect 19793 28595 19859 28598
rect 20294 28596 20300 28598
rect 20364 28658 20370 28660
rect 22645 28658 22711 28661
rect 20364 28656 22711 28658
rect 20364 28600 22650 28656
rect 22706 28600 22711 28656
rect 20364 28598 22711 28600
rect 20364 28596 20370 28598
rect 22645 28595 22711 28598
rect 29729 28658 29795 28661
rect 38009 28658 38075 28661
rect 29729 28656 38075 28658
rect 29729 28600 29734 28656
rect 29790 28600 38014 28656
rect 38070 28600 38075 28656
rect 29729 28598 38075 28600
rect 29729 28595 29795 28598
rect 38009 28595 38075 28598
rect 19701 28522 19767 28525
rect 20437 28522 20503 28525
rect 21817 28522 21883 28525
rect 22001 28522 22067 28525
rect 19701 28520 20362 28522
rect 19701 28464 19706 28520
rect 19762 28464 20362 28520
rect 19701 28462 20362 28464
rect 19701 28459 19767 28462
rect 20302 28386 20362 28462
rect 20437 28520 22067 28522
rect 20437 28464 20442 28520
rect 20498 28464 21822 28520
rect 21878 28464 22006 28520
rect 22062 28464 22067 28520
rect 20437 28462 22067 28464
rect 20437 28459 20503 28462
rect 21817 28459 21883 28462
rect 22001 28459 22067 28462
rect 20529 28386 20595 28389
rect 20302 28384 20595 28386
rect 20302 28328 20534 28384
rect 20590 28328 20595 28384
rect 20302 28326 20595 28328
rect 20529 28323 20595 28326
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 19885 28114 19951 28117
rect 22921 28114 22987 28117
rect 19885 28112 22987 28114
rect 19885 28056 19890 28112
rect 19946 28056 22926 28112
rect 22982 28056 22987 28112
rect 19885 28054 22987 28056
rect 19885 28051 19951 28054
rect 22921 28051 22987 28054
rect 19517 27978 19583 27981
rect 20897 27978 20963 27981
rect 19517 27976 20963 27978
rect 19517 27920 19522 27976
rect 19578 27920 20902 27976
rect 20958 27920 20963 27976
rect 19517 27918 20963 27920
rect 19517 27915 19583 27918
rect 20897 27915 20963 27918
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 19333 27706 19399 27709
rect 24301 27706 24367 27709
rect 19333 27704 24367 27706
rect 19333 27648 19338 27704
rect 19394 27648 24306 27704
rect 24362 27648 24367 27704
rect 19333 27646 24367 27648
rect 19333 27643 19399 27646
rect 24301 27643 24367 27646
rect 20713 27570 20779 27573
rect 21357 27570 21423 27573
rect 20713 27568 21423 27570
rect 20713 27512 20718 27568
rect 20774 27512 21362 27568
rect 21418 27512 21423 27568
rect 20713 27510 21423 27512
rect 20713 27507 20779 27510
rect 21357 27507 21423 27510
rect 19333 27434 19399 27437
rect 19885 27434 19951 27437
rect 19333 27432 19951 27434
rect 19333 27376 19338 27432
rect 19394 27376 19890 27432
rect 19946 27376 19951 27432
rect 19333 27374 19951 27376
rect 19333 27371 19399 27374
rect 19885 27371 19951 27374
rect 23565 27434 23631 27437
rect 28257 27434 28323 27437
rect 23565 27432 28323 27434
rect 23565 27376 23570 27432
rect 23626 27376 28262 27432
rect 28318 27376 28323 27432
rect 23565 27374 28323 27376
rect 23565 27371 23631 27374
rect 28257 27371 28323 27374
rect 27654 27236 27660 27300
rect 27724 27298 27730 27300
rect 27797 27298 27863 27301
rect 28349 27298 28415 27301
rect 27724 27296 28415 27298
rect 27724 27240 27802 27296
rect 27858 27240 28354 27296
rect 28410 27240 28415 27296
rect 27724 27238 28415 27240
rect 27724 27236 27730 27238
rect 27797 27235 27863 27238
rect 28349 27235 28415 27238
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 13169 27162 13235 27165
rect 17217 27162 17283 27165
rect 13169 27160 17283 27162
rect 13169 27104 13174 27160
rect 13230 27104 17222 27160
rect 17278 27104 17283 27160
rect 13169 27102 17283 27104
rect 13169 27099 13235 27102
rect 17217 27099 17283 27102
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 13353 25802 13419 25805
rect 13486 25802 13492 25804
rect 13353 25800 13492 25802
rect 13353 25744 13358 25800
rect 13414 25744 13492 25800
rect 13353 25742 13492 25744
rect 13353 25739 13419 25742
rect 13486 25740 13492 25742
rect 13556 25740 13562 25804
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 19701 25394 19767 25397
rect 21173 25394 21239 25397
rect 19701 25392 21239 25394
rect 19701 25336 19706 25392
rect 19762 25336 21178 25392
rect 21234 25336 21239 25392
rect 19701 25334 21239 25336
rect 19701 25331 19767 25334
rect 21173 25331 21239 25334
rect 27705 25260 27771 25261
rect 27654 25196 27660 25260
rect 27724 25258 27771 25260
rect 27724 25256 27816 25258
rect 27766 25200 27816 25256
rect 27724 25198 27816 25200
rect 27724 25196 27771 25198
rect 27705 25195 27771 25196
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 19517 24306 19583 24309
rect 20437 24306 20503 24309
rect 19517 24304 20503 24306
rect 19517 24248 19522 24304
rect 19578 24248 20442 24304
rect 20498 24248 20503 24304
rect 19517 24246 20503 24248
rect 19517 24243 19583 24246
rect 20437 24243 20503 24246
rect 19333 24170 19399 24173
rect 20621 24170 20687 24173
rect 25681 24170 25747 24173
rect 19333 24168 25747 24170
rect 19333 24112 19338 24168
rect 19394 24112 20626 24168
rect 20682 24112 25686 24168
rect 25742 24112 25747 24168
rect 19333 24110 25747 24112
rect 19333 24107 19399 24110
rect 20621 24107 20687 24110
rect 25681 24107 25747 24110
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 22001 23898 22067 23901
rect 24669 23898 24735 23901
rect 22001 23896 24735 23898
rect 22001 23840 22006 23896
rect 22062 23840 24674 23896
rect 24730 23840 24735 23896
rect 22001 23838 24735 23840
rect 22001 23835 22067 23838
rect 24669 23835 24735 23838
rect 19333 23762 19399 23765
rect 19517 23762 19583 23765
rect 19333 23760 19583 23762
rect 19333 23704 19338 23760
rect 19394 23704 19522 23760
rect 19578 23704 19583 23760
rect 19333 23702 19583 23704
rect 19333 23699 19399 23702
rect 19517 23699 19583 23702
rect 13905 23626 13971 23629
rect 14273 23626 14339 23629
rect 19149 23626 19215 23629
rect 13905 23624 19215 23626
rect 13905 23568 13910 23624
rect 13966 23568 14278 23624
rect 14334 23568 19154 23624
rect 19210 23568 19215 23624
rect 13905 23566 19215 23568
rect 13905 23563 13971 23566
rect 14273 23563 14339 23566
rect 19149 23563 19215 23566
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 20253 23220 20319 23221
rect 20253 23218 20300 23220
rect 20208 23216 20300 23218
rect 20208 23160 20258 23216
rect 20208 23158 20300 23160
rect 20253 23156 20300 23158
rect 20364 23156 20370 23220
rect 20253 23155 20319 23156
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 28073 22538 28139 22541
rect 28349 22538 28415 22541
rect 28073 22536 28415 22538
rect 28073 22480 28078 22536
rect 28134 22480 28354 22536
rect 28410 22480 28415 22536
rect 28073 22478 28415 22480
rect 28073 22475 28139 22478
rect 28349 22475 28415 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 28809 22132 28875 22133
rect 28758 22130 28764 22132
rect 28718 22070 28764 22130
rect 28828 22128 28875 22132
rect 28870 22072 28875 22128
rect 28758 22068 28764 22070
rect 28828 22068 28875 22072
rect 28809 22067 28875 22068
rect 23657 21994 23723 21997
rect 28809 21994 28875 21997
rect 23657 21992 28875 21994
rect 23657 21936 23662 21992
rect 23718 21936 28814 21992
rect 28870 21936 28875 21992
rect 23657 21934 28875 21936
rect 23657 21931 23723 21934
rect 28809 21931 28875 21934
rect 22737 21858 22803 21861
rect 25129 21858 25195 21861
rect 26141 21858 26207 21861
rect 22737 21856 26207 21858
rect 22737 21800 22742 21856
rect 22798 21800 25134 21856
rect 25190 21800 26146 21856
rect 26202 21800 26207 21856
rect 22737 21798 26207 21800
rect 22737 21795 22803 21798
rect 25129 21795 25195 21798
rect 26141 21795 26207 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 27705 21722 27771 21725
rect 27889 21722 27955 21725
rect 27705 21720 27955 21722
rect 27705 21664 27710 21720
rect 27766 21664 27894 21720
rect 27950 21664 27955 21720
rect 27705 21662 27955 21664
rect 27705 21659 27771 21662
rect 27889 21659 27955 21662
rect 14917 21586 14983 21589
rect 16481 21586 16547 21589
rect 27705 21588 27771 21589
rect 14917 21584 16547 21586
rect 14917 21528 14922 21584
rect 14978 21528 16486 21584
rect 16542 21528 16547 21584
rect 14917 21526 16547 21528
rect 14917 21523 14983 21526
rect 16481 21523 16547 21526
rect 27654 21524 27660 21588
rect 27724 21586 27771 21588
rect 27889 21586 27955 21589
rect 27724 21584 27955 21586
rect 27766 21528 27894 21584
rect 27950 21528 27955 21584
rect 27724 21526 27955 21528
rect 27724 21524 27771 21526
rect 27705 21523 27771 21524
rect 27889 21523 27955 21526
rect 29545 21586 29611 21589
rect 30465 21586 30531 21589
rect 29545 21584 30531 21586
rect 29545 21528 29550 21584
rect 29606 21528 30470 21584
rect 30526 21528 30531 21584
rect 29545 21526 30531 21528
rect 29545 21523 29611 21526
rect 30465 21523 30531 21526
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 25681 20906 25747 20909
rect 28073 20906 28139 20909
rect 25681 20904 28139 20906
rect 25681 20848 25686 20904
rect 25742 20848 28078 20904
rect 28134 20848 28139 20904
rect 25681 20846 28139 20848
rect 25681 20843 25747 20846
rect 28073 20843 28139 20846
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 28073 20634 28139 20637
rect 28901 20634 28967 20637
rect 28073 20632 28967 20634
rect 28073 20576 28078 20632
rect 28134 20576 28906 20632
rect 28962 20576 28967 20632
rect 28073 20574 28967 20576
rect 28073 20571 28139 20574
rect 28901 20571 28967 20574
rect 14917 20498 14983 20501
rect 16062 20498 16068 20500
rect 14917 20496 16068 20498
rect 14917 20440 14922 20496
rect 14978 20440 16068 20496
rect 14917 20438 16068 20440
rect 14917 20435 14983 20438
rect 16062 20436 16068 20438
rect 16132 20436 16138 20500
rect 20069 20498 20135 20501
rect 21357 20498 21423 20501
rect 20069 20496 21423 20498
rect 20069 20440 20074 20496
rect 20130 20440 21362 20496
rect 21418 20440 21423 20496
rect 20069 20438 21423 20440
rect 20069 20435 20135 20438
rect 21357 20435 21423 20438
rect 25405 20498 25471 20501
rect 27429 20498 27495 20501
rect 25405 20496 27495 20498
rect 25405 20440 25410 20496
rect 25466 20440 27434 20496
rect 27490 20440 27495 20496
rect 25405 20438 27495 20440
rect 25405 20435 25471 20438
rect 27429 20435 27495 20438
rect 28441 20498 28507 20501
rect 28901 20498 28967 20501
rect 28441 20496 28967 20498
rect 28441 20440 28446 20496
rect 28502 20440 28906 20496
rect 28962 20440 28967 20496
rect 28441 20438 28967 20440
rect 28441 20435 28507 20438
rect 28901 20435 28967 20438
rect 15285 20362 15351 20365
rect 15561 20362 15627 20365
rect 15285 20360 15627 20362
rect 15285 20304 15290 20360
rect 15346 20304 15566 20360
rect 15622 20304 15627 20360
rect 15285 20302 15627 20304
rect 15285 20299 15351 20302
rect 15561 20299 15627 20302
rect 29085 20362 29151 20365
rect 29085 20360 29194 20362
rect 29085 20304 29090 20360
rect 29146 20304 29194 20360
rect 29085 20299 29194 20304
rect 29134 20229 29194 20299
rect 29085 20224 29194 20229
rect 29085 20168 29090 20224
rect 29146 20168 29194 20224
rect 29085 20166 29194 20168
rect 29085 20163 29151 20166
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 20437 20092 20503 20093
rect 28717 20092 28783 20093
rect 20437 20090 20484 20092
rect 20392 20088 20484 20090
rect 20392 20032 20442 20088
rect 20392 20030 20484 20032
rect 20437 20028 20484 20030
rect 20548 20028 20554 20092
rect 28717 20090 28764 20092
rect 28672 20088 28764 20090
rect 28672 20032 28722 20088
rect 28672 20030 28764 20032
rect 28717 20028 28764 20030
rect 28828 20028 28834 20092
rect 20437 20027 20503 20028
rect 28717 20027 28783 20028
rect 27337 19818 27403 19821
rect 28349 19818 28415 19821
rect 27337 19816 28415 19818
rect 27337 19760 27342 19816
rect 27398 19760 28354 19816
rect 28410 19760 28415 19816
rect 27337 19758 28415 19760
rect 27337 19755 27403 19758
rect 28349 19755 28415 19758
rect 24761 19682 24827 19685
rect 28441 19682 28507 19685
rect 24761 19680 28507 19682
rect 24761 19624 24766 19680
rect 24822 19624 28446 19680
rect 28502 19624 28507 19680
rect 24761 19622 28507 19624
rect 24761 19619 24827 19622
rect 28441 19619 28507 19622
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 19977 19002 20043 19005
rect 20110 19002 20116 19004
rect 19977 19000 20116 19002
rect 19977 18944 19982 19000
rect 20038 18944 20116 19000
rect 19977 18942 20116 18944
rect 19977 18939 20043 18942
rect 20110 18940 20116 18942
rect 20180 18940 20186 19004
rect 19057 18866 19123 18869
rect 18462 18864 19123 18866
rect 18462 18808 19062 18864
rect 19118 18808 19123 18864
rect 18462 18806 19123 18808
rect 18321 18594 18387 18597
rect 18462 18594 18522 18806
rect 19057 18803 19123 18806
rect 18873 18730 18939 18733
rect 18873 18728 19074 18730
rect 18873 18672 18878 18728
rect 18934 18672 19074 18728
rect 18873 18670 19074 18672
rect 18873 18667 18939 18670
rect 18321 18592 18522 18594
rect 18321 18536 18326 18592
rect 18382 18536 18522 18592
rect 18321 18534 18522 18536
rect 18321 18531 18387 18534
rect 19014 18461 19074 18670
rect 19374 18668 19380 18732
rect 19444 18730 19450 18732
rect 19517 18730 19583 18733
rect 19444 18728 19583 18730
rect 19444 18672 19522 18728
rect 19578 18672 19583 18728
rect 19444 18670 19583 18672
rect 19444 18668 19450 18670
rect 19517 18667 19583 18670
rect 20069 18594 20135 18597
rect 20294 18594 20300 18596
rect 20069 18592 20300 18594
rect 20069 18536 20074 18592
rect 20130 18536 20300 18592
rect 20069 18534 20300 18536
rect 20069 18531 20135 18534
rect 20294 18532 20300 18534
rect 20364 18532 20370 18596
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 18965 18456 19074 18461
rect 18965 18400 18970 18456
rect 19026 18400 19074 18456
rect 18965 18398 19074 18400
rect 20805 18458 20871 18461
rect 20805 18456 20914 18458
rect 20805 18400 20810 18456
rect 20866 18400 20914 18456
rect 18965 18395 19031 18398
rect 20805 18395 20914 18400
rect 17585 18186 17651 18189
rect 18597 18186 18663 18189
rect 20713 18186 20779 18189
rect 17585 18184 18663 18186
rect 17585 18128 17590 18184
rect 17646 18128 18602 18184
rect 18658 18128 18663 18184
rect 17585 18126 18663 18128
rect 17585 18123 17651 18126
rect 18597 18123 18663 18126
rect 20486 18184 20779 18186
rect 20486 18128 20718 18184
rect 20774 18128 20779 18184
rect 20486 18126 20779 18128
rect 12893 18052 12959 18053
rect 12893 18048 12940 18052
rect 13004 18050 13010 18052
rect 19977 18050 20043 18053
rect 20110 18050 20116 18052
rect 12893 17992 12898 18048
rect 12893 17988 12940 17992
rect 13004 17990 13050 18050
rect 19977 18048 20116 18050
rect 19977 17992 19982 18048
rect 20038 17992 20116 18048
rect 19977 17990 20116 17992
rect 13004 17988 13010 17990
rect 12893 17987 12959 17988
rect 19977 17987 20043 17990
rect 20110 17988 20116 17990
rect 20180 17988 20186 18052
rect 20345 18050 20411 18053
rect 20486 18050 20546 18126
rect 20713 18123 20779 18126
rect 20345 18048 20546 18050
rect 20345 17992 20350 18048
rect 20406 17992 20546 18048
rect 20345 17990 20546 17992
rect 20713 18050 20779 18053
rect 20854 18050 20914 18395
rect 21081 18322 21147 18325
rect 21265 18322 21331 18325
rect 21081 18320 21331 18322
rect 21081 18264 21086 18320
rect 21142 18264 21270 18320
rect 21326 18264 21331 18320
rect 21081 18262 21331 18264
rect 21081 18259 21147 18262
rect 21265 18259 21331 18262
rect 34973 18186 35039 18189
rect 35750 18186 35756 18188
rect 34973 18184 35756 18186
rect 34973 18128 34978 18184
rect 35034 18128 35756 18184
rect 34973 18126 35756 18128
rect 34973 18123 35039 18126
rect 35750 18124 35756 18126
rect 35820 18124 35826 18188
rect 20713 18048 20914 18050
rect 20713 17992 20718 18048
rect 20774 17992 20914 18048
rect 20713 17990 20914 17992
rect 20345 17987 20411 17990
rect 20713 17987 20779 17990
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 19885 17914 19951 17917
rect 20805 17914 20871 17917
rect 19885 17912 20871 17914
rect 19885 17856 19890 17912
rect 19946 17856 20810 17912
rect 20866 17856 20871 17912
rect 19885 17854 20871 17856
rect 19885 17851 19951 17854
rect 20805 17851 20871 17854
rect 19701 17778 19767 17781
rect 24669 17778 24735 17781
rect 19701 17776 24735 17778
rect 19701 17720 19706 17776
rect 19762 17720 24674 17776
rect 24730 17720 24735 17776
rect 19701 17718 24735 17720
rect 19701 17715 19767 17718
rect 24669 17715 24735 17718
rect 9397 17508 9463 17509
rect 9397 17506 9444 17508
rect 9352 17504 9444 17506
rect 9352 17448 9402 17504
rect 9352 17446 9444 17448
rect 9397 17444 9444 17446
rect 9508 17444 9514 17508
rect 9397 17443 9463 17444
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 19517 17234 19583 17237
rect 20161 17234 20227 17237
rect 20713 17234 20779 17237
rect 19517 17232 20779 17234
rect 19517 17176 19522 17232
rect 19578 17176 20166 17232
rect 20222 17176 20718 17232
rect 20774 17176 20779 17232
rect 19517 17174 20779 17176
rect 19517 17171 19583 17174
rect 20161 17171 20227 17174
rect 20713 17171 20779 17174
rect 20069 17098 20135 17101
rect 23289 17098 23355 17101
rect 20069 17096 23355 17098
rect 20069 17040 20074 17096
rect 20130 17040 23294 17096
rect 23350 17040 23355 17096
rect 20069 17038 23355 17040
rect 20069 17035 20135 17038
rect 23289 17035 23355 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 11329 16690 11395 16693
rect 15285 16690 15351 16693
rect 16205 16690 16271 16693
rect 11329 16688 16271 16690
rect 11329 16632 11334 16688
rect 11390 16632 15290 16688
rect 15346 16632 16210 16688
rect 16266 16632 16271 16688
rect 11329 16630 16271 16632
rect 11329 16627 11395 16630
rect 15285 16627 15351 16630
rect 16205 16627 16271 16630
rect 31661 16690 31727 16693
rect 36445 16690 36511 16693
rect 31661 16688 36511 16690
rect 31661 16632 31666 16688
rect 31722 16632 36450 16688
rect 36506 16632 36511 16688
rect 31661 16630 36511 16632
rect 31661 16627 31727 16630
rect 36445 16627 36511 16630
rect 17585 16554 17651 16557
rect 17718 16554 17724 16556
rect 17585 16552 17724 16554
rect 17585 16496 17590 16552
rect 17646 16496 17724 16552
rect 17585 16494 17724 16496
rect 17585 16491 17651 16494
rect 17718 16492 17724 16494
rect 17788 16492 17794 16556
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 5257 15874 5323 15877
rect 7281 15874 7347 15877
rect 5257 15872 7347 15874
rect 5257 15816 5262 15872
rect 5318 15816 7286 15872
rect 7342 15816 7347 15872
rect 5257 15814 7347 15816
rect 5257 15811 5323 15814
rect 7281 15811 7347 15814
rect 32305 15874 32371 15877
rect 33685 15874 33751 15877
rect 32305 15872 33751 15874
rect 32305 15816 32310 15872
rect 32366 15816 33690 15872
rect 33746 15816 33751 15872
rect 32305 15814 33751 15816
rect 32305 15811 32371 15814
rect 33685 15811 33751 15814
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 30833 15602 30899 15605
rect 33869 15602 33935 15605
rect 30833 15600 33935 15602
rect 30833 15544 30838 15600
rect 30894 15544 33874 15600
rect 33930 15544 33935 15600
rect 30833 15542 33935 15544
rect 30833 15539 30899 15542
rect 33869 15539 33935 15542
rect 19374 15404 19380 15468
rect 19444 15466 19450 15468
rect 19701 15466 19767 15469
rect 19444 15464 19767 15466
rect 19444 15408 19706 15464
rect 19762 15408 19767 15464
rect 19444 15406 19767 15408
rect 19444 15404 19450 15406
rect 19701 15403 19767 15406
rect 20437 15468 20503 15469
rect 20437 15464 20484 15468
rect 20548 15466 20554 15468
rect 20437 15408 20442 15464
rect 20437 15404 20484 15408
rect 20548 15406 20594 15466
rect 20548 15404 20554 15406
rect 20437 15403 20503 15404
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 20161 15194 20227 15197
rect 20294 15194 20300 15196
rect 20161 15192 20300 15194
rect 20161 15136 20166 15192
rect 20222 15136 20300 15192
rect 20161 15134 20300 15136
rect 20161 15131 20227 15134
rect 20294 15132 20300 15134
rect 20364 15132 20370 15196
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 16481 14514 16547 14517
rect 18321 14514 18387 14517
rect 16481 14512 18387 14514
rect 16481 14456 16486 14512
rect 16542 14456 18326 14512
rect 18382 14456 18387 14512
rect 16481 14454 18387 14456
rect 16481 14451 16547 14454
rect 18321 14451 18387 14454
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 12801 12746 12867 12749
rect 14273 12746 14339 12749
rect 12801 12744 14339 12746
rect 12801 12688 12806 12744
rect 12862 12688 14278 12744
rect 14334 12688 14339 12744
rect 12801 12686 14339 12688
rect 12801 12683 12867 12686
rect 14273 12683 14339 12686
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 19374 12412 19380 12476
rect 19444 12474 19450 12476
rect 19793 12474 19859 12477
rect 19444 12472 19859 12474
rect 19444 12416 19798 12472
rect 19854 12416 19859 12472
rect 19444 12414 19859 12416
rect 19444 12412 19450 12414
rect 19793 12411 19859 12414
rect 14549 12338 14615 12341
rect 15009 12338 15075 12341
rect 18873 12338 18939 12341
rect 14549 12336 18939 12338
rect 14549 12280 14554 12336
rect 14610 12280 15014 12336
rect 15070 12280 18878 12336
rect 18934 12280 18939 12336
rect 14549 12278 18939 12280
rect 14549 12275 14615 12278
rect 15009 12275 15075 12278
rect 18873 12275 18939 12278
rect 20161 12202 20227 12205
rect 20621 12202 20687 12205
rect 20161 12200 20687 12202
rect 20161 12144 20166 12200
rect 20222 12144 20626 12200
rect 20682 12144 20687 12200
rect 20161 12142 20687 12144
rect 20161 12139 20227 12142
rect 20621 12139 20687 12142
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 26233 9618 26299 9621
rect 27521 9618 27587 9621
rect 26233 9616 27587 9618
rect 26233 9560 26238 9616
rect 26294 9560 27526 9616
rect 27582 9560 27587 9616
rect 26233 9558 27587 9560
rect 26233 9555 26299 9558
rect 27521 9555 27587 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 21265 8530 21331 8533
rect 22185 8530 22251 8533
rect 21265 8528 22251 8530
rect 21265 8472 21270 8528
rect 21326 8472 22190 8528
rect 22246 8472 22251 8528
rect 21265 8470 22251 8472
rect 21265 8467 21331 8470
rect 22185 8467 22251 8470
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 8201 8122 8267 8125
rect 13486 8122 13492 8124
rect 8201 8120 13492 8122
rect 8201 8064 8206 8120
rect 8262 8064 13492 8120
rect 8201 8062 13492 8064
rect 8201 8059 8267 8062
rect 13486 8060 13492 8062
rect 13556 8060 13562 8124
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 18597 6898 18663 6901
rect 24945 6898 25011 6901
rect 18597 6896 25011 6898
rect 18597 6840 18602 6896
rect 18658 6840 24950 6896
rect 25006 6840 25011 6896
rect 18597 6838 25011 6840
rect 18597 6835 18663 6838
rect 24945 6835 25011 6838
rect 11145 6762 11211 6765
rect 12893 6762 12959 6765
rect 11145 6760 12959 6762
rect 11145 6704 11150 6760
rect 11206 6704 12898 6760
rect 12954 6704 12959 6760
rect 11145 6702 12959 6704
rect 11145 6699 11211 6702
rect 12893 6699 12959 6702
rect 19517 6762 19583 6765
rect 21081 6762 21147 6765
rect 19517 6760 21147 6762
rect 19517 6704 19522 6760
rect 19578 6704 21086 6760
rect 21142 6704 21147 6760
rect 19517 6702 21147 6704
rect 19517 6699 19583 6702
rect 21081 6699 21147 6702
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 29453 5130 29519 5133
rect 35709 5130 35775 5133
rect 29453 5128 35775 5130
rect 29453 5072 29458 5128
rect 29514 5072 35714 5128
rect 35770 5072 35775 5128
rect 29453 5070 35775 5072
rect 29453 5067 29519 5070
rect 35709 5067 35775 5070
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 20805 4858 20871 4861
rect 22001 4858 22067 4861
rect 20805 4856 22067 4858
rect 20805 4800 20810 4856
rect 20866 4800 22006 4856
rect 22062 4800 22067 4856
rect 20805 4798 22067 4800
rect 20805 4795 20871 4798
rect 22001 4795 22067 4798
rect 19701 4722 19767 4725
rect 21725 4722 21791 4725
rect 23933 4722 23999 4725
rect 19701 4720 23999 4722
rect 19701 4664 19706 4720
rect 19762 4664 21730 4720
rect 21786 4664 23938 4720
rect 23994 4664 23999 4720
rect 19701 4662 23999 4664
rect 19701 4659 19767 4662
rect 21725 4659 21791 4662
rect 23933 4659 23999 4662
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 14641 4314 14707 4317
rect 17033 4314 17099 4317
rect 14641 4312 17099 4314
rect 14641 4256 14646 4312
rect 14702 4256 17038 4312
rect 17094 4256 17099 4312
rect 14641 4254 17099 4256
rect 14641 4251 14707 4254
rect 17033 4251 17099 4254
rect 12934 3980 12940 4044
rect 13004 4042 13010 4044
rect 15193 4042 15259 4045
rect 13004 4040 15259 4042
rect 13004 3984 15198 4040
rect 15254 3984 15259 4040
rect 13004 3982 15259 3984
rect 13004 3980 13010 3982
rect 15193 3979 15259 3982
rect 30373 4042 30439 4045
rect 34789 4042 34855 4045
rect 30373 4040 34855 4042
rect 30373 3984 30378 4040
rect 30434 3984 34794 4040
rect 34850 3984 34855 4040
rect 30373 3982 34855 3984
rect 30373 3979 30439 3982
rect 34789 3979 34855 3982
rect 35709 4044 35775 4045
rect 35709 4040 35756 4044
rect 35820 4042 35826 4044
rect 35709 3984 35714 4040
rect 35709 3980 35756 3984
rect 35820 3982 35866 4042
rect 35820 3980 35826 3982
rect 35709 3979 35775 3980
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 27521 3770 27587 3773
rect 31109 3770 31175 3773
rect 27521 3768 31175 3770
rect 27521 3712 27526 3768
rect 27582 3712 31114 3768
rect 31170 3712 31175 3768
rect 27521 3710 31175 3712
rect 27521 3707 27587 3710
rect 31109 3707 31175 3710
rect 31293 3770 31359 3773
rect 31661 3770 31727 3773
rect 31293 3768 31727 3770
rect 31293 3712 31298 3768
rect 31354 3712 31666 3768
rect 31722 3712 31727 3768
rect 31293 3710 31727 3712
rect 31293 3707 31359 3710
rect 31661 3707 31727 3710
rect 11513 3634 11579 3637
rect 9630 3632 11579 3634
rect 9630 3603 11518 3632
rect 9627 3598 11518 3603
rect 9627 3542 9632 3598
rect 9688 3576 11518 3598
rect 11574 3576 11579 3632
rect 9688 3574 11579 3576
rect 9688 3542 9693 3574
rect 11513 3571 11579 3574
rect 28441 3634 28507 3637
rect 36537 3634 36603 3637
rect 28441 3632 36603 3634
rect 28441 3576 28446 3632
rect 28502 3576 36542 3632
rect 36598 3576 36603 3632
rect 28441 3574 36603 3576
rect 28441 3571 28507 3574
rect 36537 3571 36603 3574
rect 9627 3537 9693 3542
rect 9765 3498 9831 3501
rect 10685 3498 10751 3501
rect 9765 3496 10751 3498
rect 9765 3440 9770 3496
rect 9826 3440 10690 3496
rect 10746 3440 10751 3496
rect 9765 3438 10751 3440
rect 9765 3435 9831 3438
rect 10685 3435 10751 3438
rect 19885 3498 19951 3501
rect 28809 3498 28875 3501
rect 19885 3496 28875 3498
rect 19885 3440 19890 3496
rect 19946 3440 28814 3496
rect 28870 3440 28875 3496
rect 19885 3438 28875 3440
rect 19885 3435 19951 3438
rect 28809 3435 28875 3438
rect 31109 3498 31175 3501
rect 36905 3498 36971 3501
rect 31109 3496 36971 3498
rect 31109 3440 31114 3496
rect 31170 3440 36910 3496
rect 36966 3440 36971 3496
rect 31109 3438 36971 3440
rect 31109 3435 31175 3438
rect 36905 3435 36971 3438
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 1945 2546 2011 2549
rect 9438 2546 9444 2548
rect 1945 2544 9444 2546
rect 1945 2488 1950 2544
rect 2006 2488 9444 2544
rect 1945 2486 9444 2488
rect 1945 2483 2011 2486
rect 9438 2484 9444 2486
rect 9508 2484 9514 2548
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 16068 37360 16132 37364
rect 16068 37304 16082 37360
rect 16082 37304 16132 37360
rect 16068 37300 16132 37304
rect 17724 37360 17788 37364
rect 17724 37304 17738 37360
rect 17738 37304 17788 37360
rect 17724 37300 17788 37304
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 20116 34580 20180 34644
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 20116 29820 20180 29884
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 20300 28596 20364 28660
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 27660 27236 27724 27300
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 13492 25740 13556 25804
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 27660 25256 27724 25260
rect 27660 25200 27710 25256
rect 27710 25200 27724 25256
rect 27660 25196 27724 25200
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 20300 23216 20364 23220
rect 20300 23160 20314 23216
rect 20314 23160 20364 23216
rect 20300 23156 20364 23160
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 28764 22128 28828 22132
rect 28764 22072 28814 22128
rect 28814 22072 28828 22128
rect 28764 22068 28828 22072
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 27660 21584 27724 21588
rect 27660 21528 27710 21584
rect 27710 21528 27724 21584
rect 27660 21524 27724 21528
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 16068 20436 16132 20500
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 20484 20088 20548 20092
rect 20484 20032 20498 20088
rect 20498 20032 20548 20088
rect 20484 20028 20548 20032
rect 28764 20088 28828 20092
rect 28764 20032 28778 20088
rect 28778 20032 28828 20088
rect 28764 20028 28828 20032
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 20116 18940 20180 19004
rect 19380 18668 19444 18732
rect 20300 18532 20364 18596
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 12940 18048 13004 18052
rect 12940 17992 12954 18048
rect 12954 17992 13004 18048
rect 12940 17988 13004 17992
rect 20116 17988 20180 18052
rect 35756 18124 35820 18188
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 9444 17504 9508 17508
rect 9444 17448 9458 17504
rect 9458 17448 9508 17504
rect 9444 17444 9508 17448
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 17724 16492 17788 16556
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19380 15404 19444 15468
rect 20484 15464 20548 15468
rect 20484 15408 20498 15464
rect 20498 15408 20548 15464
rect 20484 15404 20548 15408
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 20300 15132 20364 15196
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19380 12412 19444 12476
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 13492 8060 13556 8124
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 12940 3980 13004 4044
rect 35756 4040 35820 4044
rect 35756 3984 35770 4040
rect 35770 3984 35820 4040
rect 35756 3980 35820 3984
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 9444 2484 9508 2548
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 16067 37364 16133 37365
rect 16067 37300 16068 37364
rect 16132 37300 16133 37364
rect 16067 37299 16133 37300
rect 17723 37364 17789 37365
rect 17723 37300 17724 37364
rect 17788 37300 17789 37364
rect 17723 37299 17789 37300
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 13491 25804 13557 25805
rect 13491 25740 13492 25804
rect 13556 25740 13557 25804
rect 13491 25739 13557 25740
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 12939 18052 13005 18053
rect 12939 17988 12940 18052
rect 13004 17988 13005 18052
rect 12939 17987 13005 17988
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 9443 17508 9509 17509
rect 9443 17444 9444 17508
rect 9508 17444 9509 17508
rect 9443 17443 9509 17444
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 9446 2549 9506 17443
rect 12942 4045 13002 17987
rect 13494 8125 13554 25739
rect 16070 20501 16130 37299
rect 16067 20500 16133 20501
rect 16067 20436 16068 20500
rect 16132 20436 16133 20500
rect 16067 20435 16133 20436
rect 17726 16557 17786 37299
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 20115 34644 20181 34645
rect 20115 34580 20116 34644
rect 20180 34580 20181 34644
rect 20115 34579 20181 34580
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 20118 29885 20178 34579
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 20115 29884 20181 29885
rect 20115 29820 20116 29884
rect 20180 29820 20181 29884
rect 20115 29819 20181 29820
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 20299 28660 20365 28661
rect 20299 28596 20300 28660
rect 20364 28596 20365 28660
rect 20299 28595 20365 28596
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 20302 23221 20362 28595
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 27659 27300 27725 27301
rect 27659 27236 27660 27300
rect 27724 27236 27725 27300
rect 27659 27235 27725 27236
rect 27662 25261 27722 27235
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 27659 25260 27725 25261
rect 27659 25196 27660 25260
rect 27724 25196 27725 25260
rect 27659 25195 27725 25196
rect 20299 23220 20365 23221
rect 20299 23156 20300 23220
rect 20364 23156 20365 23220
rect 20299 23155 20365 23156
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 27662 21589 27722 25195
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 28763 22132 28829 22133
rect 28763 22068 28764 22132
rect 28828 22068 28829 22132
rect 28763 22067 28829 22068
rect 27659 21588 27725 21589
rect 27659 21524 27660 21588
rect 27724 21524 27725 21588
rect 27659 21523 27725 21524
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 28766 20093 28826 22067
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 20483 20092 20549 20093
rect 20483 20028 20484 20092
rect 20548 20028 20549 20092
rect 20483 20027 20549 20028
rect 28763 20092 28829 20093
rect 28763 20028 28764 20092
rect 28828 20028 28829 20092
rect 28763 20027 28829 20028
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19379 18732 19445 18733
rect 19379 18668 19380 18732
rect 19444 18668 19445 18732
rect 19379 18667 19445 18668
rect 17723 16556 17789 16557
rect 17723 16492 17724 16556
rect 17788 16492 17789 16556
rect 17723 16491 17789 16492
rect 19382 15469 19442 18667
rect 19568 18528 19888 19552
rect 20115 19004 20181 19005
rect 20115 18940 20116 19004
rect 20180 18940 20181 19004
rect 20115 18939 20181 18940
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 20118 18053 20178 18939
rect 20299 18596 20365 18597
rect 20299 18532 20300 18596
rect 20364 18532 20365 18596
rect 20299 18531 20365 18532
rect 20115 18052 20181 18053
rect 20115 17988 20116 18052
rect 20180 17988 20181 18052
rect 20115 17987 20181 17988
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19379 15468 19445 15469
rect 19379 15404 19380 15468
rect 19444 15404 19445 15468
rect 19379 15403 19445 15404
rect 19382 12477 19442 15403
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 20302 15197 20362 18531
rect 20486 15469 20546 20027
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 35755 18188 35821 18189
rect 35755 18124 35756 18188
rect 35820 18124 35821 18188
rect 35755 18123 35821 18124
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 20483 15468 20549 15469
rect 20483 15404 20484 15468
rect 20548 15404 20549 15468
rect 20483 15403 20549 15404
rect 20299 15196 20365 15197
rect 20299 15132 20300 15196
rect 20364 15132 20365 15196
rect 20299 15131 20365 15132
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19379 12476 19445 12477
rect 19379 12412 19380 12476
rect 19444 12412 19445 12476
rect 19379 12411 19445 12412
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 13491 8124 13557 8125
rect 13491 8060 13492 8124
rect 13556 8060 13557 8124
rect 13491 8059 13557 8060
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 12939 4044 13005 4045
rect 12939 3980 12940 4044
rect 13004 3980 13005 4044
rect 12939 3979 13005 3980
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 9443 2548 9509 2549
rect 9443 2484 9444 2548
rect 9508 2484 9509 2548
rect 9443 2483 9509 2484
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 35758 4045 35818 18123
rect 35755 4044 35821 4045
rect 35755 3980 35756 4044
rect 35820 3980 35821 4044
rect 35755 3979 35821 3980
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform -1 0 5244 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 12328 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform 1 0 15364 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform -1 0 19688 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform -1 0 17480 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1644511149
transform 1 0 12696 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1644511149
transform 1 0 25024 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4324 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1644511149
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67
timestamp 1644511149
transform 1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7912 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1644511149
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89
timestamp 1644511149
transform 1 0 9292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99
timestamp 1644511149
transform 1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106
timestamp 1644511149
transform 1 0 10856 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1644511149
transform 1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_135
timestamp 1644511149
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1644511149
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_150
timestamp 1644511149
transform 1 0 14904 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_158
timestamp 1644511149
transform 1 0 15640 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1644511149
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_174
timestamp 1644511149
transform 1 0 17112 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_184
timestamp 1644511149
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1644511149
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_202
timestamp 1644511149
transform 1 0 19688 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_210
timestamp 1644511149
transform 1 0 20424 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 1644511149
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1644511149
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_229
timestamp 1644511149
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_237
timestamp 1644511149
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_246
timestamp 1644511149
transform 1 0 23736 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_259
timestamp 1644511149
transform 1 0 24932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_270
timestamp 1644511149
transform 1 0 25944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1644511149
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_285
timestamp 1644511149
transform 1 0 27324 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_298
timestamp 1644511149
transform 1 0 28520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1644511149
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_317
timestamp 1644511149
transform 1 0 30268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_325
timestamp 1644511149
transform 1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1644511149
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_342
timestamp 1644511149
transform 1 0 32568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_350
timestamp 1644511149
transform 1 0 33304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_358
timestamp 1644511149
transform 1 0 34040 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_369
timestamp 1644511149
transform 1 0 35052 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_388
timestamp 1644511149
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1644511149
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_7
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_14
timestamp 1644511149
transform 1 0 2392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_18
timestamp 1644511149
transform 1 0 2760 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_25
timestamp 1644511149
transform 1 0 3404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_32
timestamp 1644511149
transform 1 0 4048 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_41
timestamp 1644511149
transform 1 0 4876 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_45
timestamp 1644511149
transform 1 0 5244 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1644511149
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_60
timestamp 1644511149
transform 1 0 6624 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_68
timestamp 1644511149
transform 1 0 7360 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_86
timestamp 1644511149
transform 1 0 9016 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_94
timestamp 1644511149
transform 1 0 9752 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_99
timestamp 1644511149
transform 1 0 10212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1644511149
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_120
timestamp 1644511149
transform 1 0 12144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_129
timestamp 1644511149
transform 1 0 12972 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_133
timestamp 1644511149
transform 1 0 13340 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_150
timestamp 1644511149
transform 1 0 14904 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_158
timestamp 1644511149
transform 1 0 15640 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1644511149
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_176
timestamp 1644511149
transform 1 0 17296 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_198
timestamp 1644511149
transform 1 0 19320 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_209
timestamp 1644511149
transform 1 0 20332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1644511149
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_233
timestamp 1644511149
transform 1 0 22540 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_240
timestamp 1644511149
transform 1 0 23184 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_251
timestamp 1644511149
transform 1 0 24196 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_259
timestamp 1644511149
transform 1 0 24932 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1644511149
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_301
timestamp 1644511149
transform 1 0 28796 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_309
timestamp 1644511149
transform 1 0 29532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_326
timestamp 1644511149
transform 1 0 31096 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1644511149
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_353
timestamp 1644511149
transform 1 0 33580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_373
timestamp 1644511149
transform 1 0 35420 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_381
timestamp 1644511149
transform 1 0 36156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1644511149
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1644511149
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_6
timestamp 1644511149
transform 1 0 1656 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_14
timestamp 1644511149
transform 1 0 2392 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_18
timestamp 1644511149
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1644511149
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1644511149
transform 1 0 5152 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_56
timestamp 1644511149
transform 1 0 6256 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_62
timestamp 1644511149
transform 1 0 6808 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_73
timestamp 1644511149
transform 1 0 7820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1644511149
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_90
timestamp 1644511149
transform 1 0 9384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_110
timestamp 1644511149
transform 1 0 11224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_130
timestamp 1644511149
transform 1 0 13064 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1644511149
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_146
timestamp 1644511149
transform 1 0 14536 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_154
timestamp 1644511149
transform 1 0 15272 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_172
timestamp 1644511149
transform 1 0 16928 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_179
timestamp 1644511149
transform 1 0 17572 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_190
timestamp 1644511149
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_201
timestamp 1644511149
transform 1 0 19596 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_221
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_228
timestamp 1644511149
transform 1 0 22080 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1644511149
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_260
timestamp 1644511149
transform 1 0 25024 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_268
timestamp 1644511149
transform 1 0 25760 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_279
timestamp 1644511149
transform 1 0 26772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_286
timestamp 1644511149
transform 1 0 27416 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_295
timestamp 1644511149
transform 1 0 28244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_302
timestamp 1644511149
transform 1 0 28888 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_318
timestamp 1644511149
transform 1 0 30360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_326
timestamp 1644511149
transform 1 0 31096 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_341
timestamp 1644511149
transform 1 0 32476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_348
timestamp 1644511149
transform 1 0 33120 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_354
timestamp 1644511149
transform 1 0 33672 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1644511149
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_372
timestamp 1644511149
transform 1 0 35328 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_380
timestamp 1644511149
transform 1 0 36064 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_384
timestamp 1644511149
transform 1 0 36432 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_397
timestamp 1644511149
transform 1 0 37628 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_403
timestamp 1644511149
transform 1 0 38180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_10
timestamp 1644511149
transform 1 0 2024 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_22
timestamp 1644511149
transform 1 0 3128 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_34
timestamp 1644511149
transform 1 0 4232 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_46
timestamp 1644511149
transform 1 0 5336 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1644511149
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_97
timestamp 1644511149
transform 1 0 10028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_106
timestamp 1644511149
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_120
timestamp 1644511149
transform 1 0 12144 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_131
timestamp 1644511149
transform 1 0 13156 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_142
timestamp 1644511149
transform 1 0 14168 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_146
timestamp 1644511149
transform 1 0 14536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_151
timestamp 1644511149
transform 1 0 14996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_172
timestamp 1644511149
transform 1 0 16928 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_188
timestamp 1644511149
transform 1 0 18400 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_200
timestamp 1644511149
transform 1 0 19504 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_206
timestamp 1644511149
transform 1 0 20056 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_211
timestamp 1644511149
transform 1 0 20516 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_218
timestamp 1644511149
transform 1 0 21160 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_241
timestamp 1644511149
transform 1 0 23276 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_247
timestamp 1644511149
transform 1 0 23828 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_252
timestamp 1644511149
transform 1 0 24288 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_266
timestamp 1644511149
transform 1 0 25576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_274
timestamp 1644511149
transform 1 0 26312 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_285
timestamp 1644511149
transform 1 0 27324 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_300
timestamp 1644511149
transform 1 0 28704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_306
timestamp 1644511149
transform 1 0 29256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_314
timestamp 1644511149
transform 1 0 29992 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_325
timestamp 1644511149
transform 1 0 31004 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_332
timestamp 1644511149
transform 1 0 31648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_340
timestamp 1644511149
transform 1 0 32384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_347
timestamp 1644511149
transform 1 0 33028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_354
timestamp 1644511149
transform 1 0 33672 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_360
timestamp 1644511149
transform 1 0 34224 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_366
timestamp 1644511149
transform 1 0 34776 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_380
timestamp 1644511149
transform 1 0 36064 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_384
timestamp 1644511149
transform 1 0 36432 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1644511149
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_401
timestamp 1644511149
transform 1 0 37996 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_89
timestamp 1644511149
transform 1 0 9292 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_102
timestamp 1644511149
transform 1 0 10488 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_110
timestamp 1644511149
transform 1 0 11224 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_114
timestamp 1644511149
transform 1 0 11592 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_118
timestamp 1644511149
transform 1 0 11960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_122
timestamp 1644511149
transform 1 0 12328 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_129
timestamp 1644511149
transform 1 0 12972 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1644511149
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_146
timestamp 1644511149
transform 1 0 14536 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_159
timestamp 1644511149
transform 1 0 15732 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_166
timestamp 1644511149
transform 1 0 16376 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_170
timestamp 1644511149
transform 1 0 16744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_187
timestamp 1644511149
transform 1 0 18308 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_200
timestamp 1644511149
transform 1 0 19504 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_207
timestamp 1644511149
transform 1 0 20148 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_215
timestamp 1644511149
transform 1 0 20884 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_220
timestamp 1644511149
transform 1 0 21344 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_229
timestamp 1644511149
transform 1 0 22172 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_237
timestamp 1644511149
transform 1 0 22908 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_258
timestamp 1644511149
transform 1 0 24840 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_267
timestamp 1644511149
transform 1 0 25668 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_280
timestamp 1644511149
transform 1 0 26864 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_287
timestamp 1644511149
transform 1 0 27508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_294
timestamp 1644511149
transform 1 0 28152 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1644511149
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_331
timestamp 1644511149
transform 1 0 31556 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_339
timestamp 1644511149
transform 1 0 32292 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_346
timestamp 1644511149
transform 1 0 32936 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_352
timestamp 1644511149
transform 1 0 33488 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_356
timestamp 1644511149
transform 1 0 33856 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_372
timestamp 1644511149
transform 1 0 35328 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_379
timestamp 1644511149
transform 1 0 35972 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_391
timestamp 1644511149
transform 1 0 37076 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_395
timestamp 1644511149
transform 1 0 37444 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_403
timestamp 1644511149
transform 1 0 38180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_89
timestamp 1644511149
transform 1 0 9292 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_94
timestamp 1644511149
transform 1 0 9752 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_102
timestamp 1644511149
transform 1 0 10488 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_106
timestamp 1644511149
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_118
timestamp 1644511149
transform 1 0 11960 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_140
timestamp 1644511149
transform 1 0 13984 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 1644511149
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_178
timestamp 1644511149
transform 1 0 17480 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_187
timestamp 1644511149
transform 1 0 18308 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_194
timestamp 1644511149
transform 1 0 18952 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_203
timestamp 1644511149
transform 1 0 19780 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_207
timestamp 1644511149
transform 1 0 20148 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_211
timestamp 1644511149
transform 1 0 20516 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_219
timestamp 1644511149
transform 1 0 21252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_228
timestamp 1644511149
transform 1 0 22080 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_238
timestamp 1644511149
transform 1 0 23000 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_258
timestamp 1644511149
transform 1 0 24840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_266
timestamp 1644511149
transform 1 0 25576 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_272
timestamp 1644511149
transform 1 0 26128 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1644511149
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_297
timestamp 1644511149
transform 1 0 28428 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_324
timestamp 1644511149
transform 1 0 30912 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_328
timestamp 1644511149
transform 1 0 31280 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_332
timestamp 1644511149
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_353
timestamp 1644511149
transform 1 0 33580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_365
timestamp 1644511149
transform 1 0 34684 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_372
timestamp 1644511149
transform 1 0 35328 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_384
timestamp 1644511149
transform 1 0 36432 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_403
timestamp 1644511149
transform 1 0 38180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_90
timestamp 1644511149
transform 1 0 9384 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_99
timestamp 1644511149
transform 1 0 10212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_108
timestamp 1644511149
transform 1 0 11040 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_119
timestamp 1644511149
transform 1 0 12052 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_125
timestamp 1644511149
transform 1 0 12604 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1644511149
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_163
timestamp 1644511149
transform 1 0 16100 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_170
timestamp 1644511149
transform 1 0 16744 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_184
timestamp 1644511149
transform 1 0 18032 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_188
timestamp 1644511149
transform 1 0 18400 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 1644511149
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_213
timestamp 1644511149
transform 1 0 20700 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_226
timestamp 1644511149
transform 1 0 21896 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_234
timestamp 1644511149
transform 1 0 22632 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_242
timestamp 1644511149
transform 1 0 23368 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_248
timestamp 1644511149
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_256
timestamp 1644511149
transform 1 0 24656 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_270
timestamp 1644511149
transform 1 0 25944 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_279
timestamp 1644511149
transform 1 0 26772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_286
timestamp 1644511149
transform 1 0 27416 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_294
timestamp 1644511149
transform 1 0 28152 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_312
timestamp 1644511149
transform 1 0 29808 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_319
timestamp 1644511149
transform 1 0 30452 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_326
timestamp 1644511149
transform 1 0 31096 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_359
timestamp 1644511149
transform 1 0 34132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_381
timestamp 1644511149
transform 1 0 36156 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_393
timestamp 1644511149
transform 1 0 37260 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_399
timestamp 1644511149
transform 1 0 37812 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_403
timestamp 1644511149
transform 1 0 38180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_75
timestamp 1644511149
transform 1 0 8004 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_95
timestamp 1644511149
transform 1 0 9844 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1644511149
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_131
timestamp 1644511149
transform 1 0 13156 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_138
timestamp 1644511149
transform 1 0 13800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_145
timestamp 1644511149
transform 1 0 14444 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_151
timestamp 1644511149
transform 1 0 14996 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_155
timestamp 1644511149
transform 1 0 15364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_174
timestamp 1644511149
transform 1 0 17112 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_196
timestamp 1644511149
transform 1 0 19136 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_204
timestamp 1644511149
transform 1 0 19872 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_210
timestamp 1644511149
transform 1 0 20424 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1644511149
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_232
timestamp 1644511149
transform 1 0 22448 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_239
timestamp 1644511149
transform 1 0 23092 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_243
timestamp 1644511149
transform 1 0 23460 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_247
timestamp 1644511149
transform 1 0 23828 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_251
timestamp 1644511149
transform 1 0 24196 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_256
timestamp 1644511149
transform 1 0 24656 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1644511149
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_289
timestamp 1644511149
transform 1 0 27692 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_296
timestamp 1644511149
transform 1 0 28336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_304
timestamp 1644511149
transform 1 0 29072 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_312
timestamp 1644511149
transform 1 0 29808 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_316
timestamp 1644511149
transform 1 0 30176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_320
timestamp 1644511149
transform 1 0 30544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_327
timestamp 1644511149
transform 1 0 31188 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_343
timestamp 1644511149
transform 1 0 32660 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_352
timestamp 1644511149
transform 1 0 33488 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_359
timestamp 1644511149
transform 1 0 34132 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_371
timestamp 1644511149
transform 1 0 35236 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_383
timestamp 1644511149
transform 1 0 36340 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_91
timestamp 1644511149
transform 1 0 9476 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_111
timestamp 1644511149
transform 1 0 11316 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_120
timestamp 1644511149
transform 1 0 12144 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_127
timestamp 1644511149
transform 1 0 12788 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1644511149
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_159
timestamp 1644511149
transform 1 0 15732 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_180
timestamp 1644511149
transform 1 0 17664 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_187
timestamp 1644511149
transform 1 0 18308 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_204
timestamp 1644511149
transform 1 0 19872 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_225
timestamp 1644511149
transform 1 0 21804 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1644511149
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_256
timestamp 1644511149
transform 1 0 24656 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_263
timestamp 1644511149
transform 1 0 25300 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_270
timestamp 1644511149
transform 1 0 25944 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_274
timestamp 1644511149
transform 1 0 26312 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_295
timestamp 1644511149
transform 1 0 28244 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_302
timestamp 1644511149
transform 1 0 28888 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_316
timestamp 1644511149
transform 1 0 30176 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_325
timestamp 1644511149
transform 1 0 31004 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_334
timestamp 1644511149
transform 1 0 31832 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_356
timestamp 1644511149
transform 1 0 33856 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_371
timestamp 1644511149
transform 1 0 35236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_383
timestamp 1644511149
transform 1 0 36340 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_395
timestamp 1644511149
transform 1 0 37444 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_82
timestamp 1644511149
transform 1 0 8648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_91
timestamp 1644511149
transform 1 0 9476 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_103
timestamp 1644511149
transform 1 0 10580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_121
timestamp 1644511149
transform 1 0 12236 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_131
timestamp 1644511149
transform 1 0 13156 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_151
timestamp 1644511149
transform 1 0 14996 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_159
timestamp 1644511149
transform 1 0 15732 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_177
timestamp 1644511149
transform 1 0 17388 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_189
timestamp 1644511149
transform 1 0 18492 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_197
timestamp 1644511149
transform 1 0 19228 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_212
timestamp 1644511149
transform 1 0 20608 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1644511149
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_234
timestamp 1644511149
transform 1 0 22632 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_242
timestamp 1644511149
transform 1 0 23368 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_257
timestamp 1644511149
transform 1 0 24748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_268
timestamp 1644511149
transform 1 0 25760 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp 1644511149
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_286
timestamp 1644511149
transform 1 0 27416 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_304
timestamp 1644511149
transform 1 0 29072 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_311
timestamp 1644511149
transform 1 0 29716 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_332
timestamp 1644511149
transform 1 0 31648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_341
timestamp 1644511149
transform 1 0 32476 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_345
timestamp 1644511149
transform 1 0 32844 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_357
timestamp 1644511149
transform 1 0 33948 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_363
timestamp 1644511149
transform 1 0 34500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_371
timestamp 1644511149
transform 1 0 35236 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_383
timestamp 1644511149
transform 1 0 36340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_61
timestamp 1644511149
transform 1 0 6716 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_79
timestamp 1644511149
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_100
timestamp 1644511149
transform 1 0 10304 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_113
timestamp 1644511149
transform 1 0 11500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_119
timestamp 1644511149
transform 1 0 12052 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_131
timestamp 1644511149
transform 1 0 13156 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_152
timestamp 1644511149
transform 1 0 15088 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_159
timestamp 1644511149
transform 1 0 15732 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_171
timestamp 1644511149
transform 1 0 16836 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_183
timestamp 1644511149
transform 1 0 17940 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1644511149
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_205
timestamp 1644511149
transform 1 0 19964 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_211
timestamp 1644511149
transform 1 0 20516 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_219
timestamp 1644511149
transform 1 0 21252 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_226
timestamp 1644511149
transform 1 0 21896 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_235
timestamp 1644511149
transform 1 0 22724 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_239
timestamp 1644511149
transform 1 0 23092 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_244
timestamp 1644511149
transform 1 0 23552 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_257
timestamp 1644511149
transform 1 0 24748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_264
timestamp 1644511149
transform 1 0 25392 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_283
timestamp 1644511149
transform 1 0 27140 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1644511149
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_329
timestamp 1644511149
transform 1 0 31372 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_337
timestamp 1644511149
transform 1 0 32108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_341
timestamp 1644511149
transform 1 0 32476 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_350
timestamp 1644511149
transform 1 0 33304 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_356
timestamp 1644511149
transform 1 0 33856 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_360
timestamp 1644511149
transform 1 0 34224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_381
timestamp 1644511149
transform 1 0 36156 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_393
timestamp 1644511149
transform 1 0 37260 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1644511149
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_72
timestamp 1644511149
transform 1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_76
timestamp 1644511149
transform 1 0 8096 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_84
timestamp 1644511149
transform 1 0 8832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1644511149
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_120
timestamp 1644511149
transform 1 0 12144 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_142
timestamp 1644511149
transform 1 0 14168 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_146
timestamp 1644511149
transform 1 0 14536 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1644511149
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_177
timestamp 1644511149
transform 1 0 17388 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_185
timestamp 1644511149
transform 1 0 18124 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_196
timestamp 1644511149
transform 1 0 19136 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_203
timestamp 1644511149
transform 1 0 19780 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_260
timestamp 1644511149
transform 1 0 25024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_268
timestamp 1644511149
transform 1 0 25760 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_272
timestamp 1644511149
transform 1 0 26128 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1644511149
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_297
timestamp 1644511149
transform 1 0 28428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_313
timestamp 1644511149
transform 1 0 29900 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_325
timestamp 1644511149
transform 1 0 31004 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_333
timestamp 1644511149
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_341
timestamp 1644511149
transform 1 0 32476 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_358
timestamp 1644511149
transform 1 0 34040 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_369
timestamp 1644511149
transform 1 0 35052 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_381
timestamp 1644511149
transform 1 0 36156 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp 1644511149
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_90
timestamp 1644511149
transform 1 0 9384 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_111
timestamp 1644511149
transform 1 0 11316 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_132
timestamp 1644511149
transform 1 0 13248 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_152
timestamp 1644511149
transform 1 0 15088 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_159
timestamp 1644511149
transform 1 0 15732 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_169
timestamp 1644511149
transform 1 0 16652 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_183
timestamp 1644511149
transform 1 0 17940 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1644511149
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_214
timestamp 1644511149
transform 1 0 20792 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_223
timestamp 1644511149
transform 1 0 21620 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_234
timestamp 1644511149
transform 1 0 22632 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1644511149
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_270
timestamp 1644511149
transform 1 0 25944 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_282
timestamp 1644511149
transform 1 0 27048 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_293
timestamp 1644511149
transform 1 0 28060 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_305
timestamp 1644511149
transform 1 0 29164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_342
timestamp 1644511149
transform 1 0 32568 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_352
timestamp 1644511149
transform 1 0 33488 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_73
timestamp 1644511149
transform 1 0 7820 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_91
timestamp 1644511149
transform 1 0 9476 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_97
timestamp 1644511149
transform 1 0 10028 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_101
timestamp 1644511149
transform 1 0 10396 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1644511149
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_119
timestamp 1644511149
transform 1 0 12052 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_127
timestamp 1644511149
transform 1 0 12788 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_134
timestamp 1644511149
transform 1 0 13432 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_146
timestamp 1644511149
transform 1 0 14536 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_154
timestamp 1644511149
transform 1 0 15272 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1644511149
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_177
timestamp 1644511149
transform 1 0 17388 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_197
timestamp 1644511149
transform 1 0 19228 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_201
timestamp 1644511149
transform 1 0 19596 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_206
timestamp 1644511149
transform 1 0 20056 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_214
timestamp 1644511149
transform 1 0 20792 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_218
timestamp 1644511149
transform 1 0 21160 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_242
timestamp 1644511149
transform 1 0 23368 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_250
timestamp 1644511149
transform 1 0 24104 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_257
timestamp 1644511149
transform 1 0 24748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_265
timestamp 1644511149
transform 1 0 25484 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_274
timestamp 1644511149
transform 1 0 26312 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_286
timestamp 1644511149
transform 1 0 27416 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_314
timestamp 1644511149
transform 1 0 29992 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_322
timestamp 1644511149
transform 1 0 30728 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_328
timestamp 1644511149
transform 1 0 31280 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_340
timestamp 1644511149
transform 1 0 32384 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_352
timestamp 1644511149
transform 1 0 33488 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_364
timestamp 1644511149
transform 1 0 34592 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_376
timestamp 1644511149
transform 1 0 35696 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_388
timestamp 1644511149
transform 1 0 36800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1644511149
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_11
timestamp 1644511149
transform 1 0 2116 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1644511149
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_88
timestamp 1644511149
transform 1 0 9200 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_100
timestamp 1644511149
transform 1 0 10304 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_104
timestamp 1644511149
transform 1 0 10672 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_111
timestamp 1644511149
transform 1 0 11316 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_123
timestamp 1644511149
transform 1 0 12420 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_129
timestamp 1644511149
transform 1 0 12972 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1644511149
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_152
timestamp 1644511149
transform 1 0 15088 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_160
timestamp 1644511149
transform 1 0 15824 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_169
timestamp 1644511149
transform 1 0 16652 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1644511149
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_228
timestamp 1644511149
transform 1 0 22080 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_240
timestamp 1644511149
transform 1 0 23184 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_261
timestamp 1644511149
transform 1 0 25116 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_282
timestamp 1644511149
transform 1 0 27048 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1644511149
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_319
timestamp 1644511149
transform 1 0 30452 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_326
timestamp 1644511149
transform 1 0 31096 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_334
timestamp 1644511149
transform 1 0 31832 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_339
timestamp 1644511149
transform 1 0 32292 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_359
timestamp 1644511149
transform 1 0 34132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_99
timestamp 1644511149
transform 1 0 10212 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1644511149
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_130
timestamp 1644511149
transform 1 0 13064 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_138
timestamp 1644511149
transform 1 0 13800 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_147
timestamp 1644511149
transform 1 0 14628 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1644511149
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_178
timestamp 1644511149
transform 1 0 17480 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_190
timestamp 1644511149
transform 1 0 18584 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_201
timestamp 1644511149
transform 1 0 19596 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1644511149
transform 1 0 20240 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1644511149
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_245
timestamp 1644511149
transform 1 0 23644 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_252
timestamp 1644511149
transform 1 0 24288 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_256
timestamp 1644511149
transform 1 0 24656 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_262
timestamp 1644511149
transform 1 0 25208 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_274
timestamp 1644511149
transform 1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_292
timestamp 1644511149
transform 1 0 27968 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_304
timestamp 1644511149
transform 1 0 29072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_311
timestamp 1644511149
transform 1 0 29716 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_319
timestamp 1644511149
transform 1 0 30452 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_326
timestamp 1644511149
transform 1 0 31096 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1644511149
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_359
timestamp 1644511149
transform 1 0 34132 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_371
timestamp 1644511149
transform 1 0 35236 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_383
timestamp 1644511149
transform 1 0 36340 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_93
timestamp 1644511149
transform 1 0 9660 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_99
timestamp 1644511149
transform 1 0 10212 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_111
timestamp 1644511149
transform 1 0 11316 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1644511149
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1644511149
transform 1 0 14812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_158
timestamp 1644511149
transform 1 0 15640 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_167
timestamp 1644511149
transform 1 0 16468 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_171
timestamp 1644511149
transform 1 0 16836 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_179
timestamp 1644511149
transform 1 0 17572 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_214
timestamp 1644511149
transform 1 0 20792 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_223
timestamp 1644511149
transform 1 0 21620 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_235
timestamp 1644511149
transform 1 0 22724 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1644511149
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_269
timestamp 1644511149
transform 1 0 25852 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_281
timestamp 1644511149
transform 1 0 26956 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_299
timestamp 1644511149
transform 1 0 28612 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_313
timestamp 1644511149
transform 1 0 29900 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_330
timestamp 1644511149
transform 1 0 31464 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_338
timestamp 1644511149
transform 1 0 32200 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_360
timestamp 1644511149
transform 1 0 34224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_73
timestamp 1644511149
transform 1 0 7820 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_77
timestamp 1644511149
transform 1 0 8188 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_89
timestamp 1644511149
transform 1 0 9292 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_101
timestamp 1644511149
transform 1 0 10396 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 1644511149
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_121
timestamp 1644511149
transform 1 0 12236 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_129
timestamp 1644511149
transform 1 0 12972 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_143
timestamp 1644511149
transform 1 0 14260 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1644511149
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_177
timestamp 1644511149
transform 1 0 17388 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_189
timestamp 1644511149
transform 1 0 18492 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_197
timestamp 1644511149
transform 1 0 19228 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_206
timestamp 1644511149
transform 1 0 20056 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_214
timestamp 1644511149
transform 1 0 20792 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1644511149
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_242
timestamp 1644511149
transform 1 0 23368 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_262
timestamp 1644511149
transform 1 0 25208 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1644511149
transform 1 0 25852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_277
timestamp 1644511149
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_284
timestamp 1644511149
transform 1 0 27232 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_301
timestamp 1644511149
transform 1 0 28796 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_313
timestamp 1644511149
transform 1 0 29900 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_325
timestamp 1644511149
transform 1 0 31004 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1644511149
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_359
timestamp 1644511149
transform 1 0 34132 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_366
timestamp 1644511149
transform 1 0 34776 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_378
timestamp 1644511149
transform 1 0 35880 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1644511149
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_61
timestamp 1644511149
transform 1 0 6716 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1644511149
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1644511149
transform 1 0 9476 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_95
timestamp 1644511149
transform 1 0 9844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_102
timestamp 1644511149
transform 1 0 10488 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_114
timestamp 1644511149
transform 1 0 11592 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_126
timestamp 1644511149
transform 1 0 12696 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1644511149
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_146
timestamp 1644511149
transform 1 0 14536 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_159
timestamp 1644511149
transform 1 0 15732 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_167
timestamp 1644511149
transform 1 0 16468 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_180
timestamp 1644511149
transform 1 0 17664 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_188
timestamp 1644511149
transform 1 0 18400 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_205
timestamp 1644511149
transform 1 0 19964 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_227
timestamp 1644511149
transform 1 0 21988 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_240
timestamp 1644511149
transform 1 0 23184 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_247
timestamp 1644511149
transform 1 0 23828 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_262
timestamp 1644511149
transform 1 0 25208 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_282
timestamp 1644511149
transform 1 0 27048 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_286
timestamp 1644511149
transform 1 0 27416 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_297
timestamp 1644511149
transform 1 0 28428 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1644511149
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_312
timestamp 1644511149
transform 1 0 29808 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_325
timestamp 1644511149
transform 1 0 31004 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_334
timestamp 1644511149
transform 1 0 31832 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_347
timestamp 1644511149
transform 1 0 33028 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_356
timestamp 1644511149
transform 1 0 33856 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_33
timestamp 1644511149
transform 1 0 4140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1644511149
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1644511149
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_65
timestamp 1644511149
transform 1 0 7084 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_84
timestamp 1644511149
transform 1 0 8832 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_92
timestamp 1644511149
transform 1 0 9568 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_96
timestamp 1644511149
transform 1 0 9936 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_102
timestamp 1644511149
transform 1 0 10488 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1644511149
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_123
timestamp 1644511149
transform 1 0 12420 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_130
timestamp 1644511149
transform 1 0 13064 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_142
timestamp 1644511149
transform 1 0 14168 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_157
timestamp 1644511149
transform 1 0 15548 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 1644511149
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1644511149
transform 1 0 17480 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_190
timestamp 1644511149
transform 1 0 18584 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_200
timestamp 1644511149
transform 1 0 19504 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_208
timestamp 1644511149
transform 1 0 20240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_215
timestamp 1644511149
transform 1 0 20884 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_248
timestamp 1644511149
transform 1 0 23920 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_260
timestamp 1644511149
transform 1 0 25024 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_272
timestamp 1644511149
transform 1 0 26128 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_298
timestamp 1644511149
transform 1 0 28520 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_341
timestamp 1644511149
transform 1 0 32476 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_347
timestamp 1644511149
transform 1 0 33028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_359
timestamp 1644511149
transform 1 0 34132 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_371
timestamp 1644511149
transform 1 0 35236 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_383
timestamp 1644511149
transform 1 0 36340 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_59
timestamp 1644511149
transform 1 0 6532 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_63
timestamp 1644511149
transform 1 0 6900 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1644511149
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_90
timestamp 1644511149
transform 1 0 9384 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_96
timestamp 1644511149
transform 1 0 9936 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_114
timestamp 1644511149
transform 1 0 11592 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_118
timestamp 1644511149
transform 1 0 11960 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1644511149
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_144
timestamp 1644511149
transform 1 0 14352 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_171
timestamp 1644511149
transform 1 0 16836 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_181
timestamp 1644511149
transform 1 0 17756 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_204
timestamp 1644511149
transform 1 0 19872 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_216
timestamp 1644511149
transform 1 0 20976 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_228
timestamp 1644511149
transform 1 0 22080 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_240
timestamp 1644511149
transform 1 0 23184 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_244
timestamp 1644511149
transform 1 0 23552 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1644511149
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_257
timestamp 1644511149
transform 1 0 24748 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_269
timestamp 1644511149
transform 1 0 25852 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_285
timestamp 1644511149
transform 1 0 27324 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_292
timestamp 1644511149
transform 1 0 27968 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_304
timestamp 1644511149
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_320
timestamp 1644511149
transform 1 0 30544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_327
timestamp 1644511149
transform 1 0 31188 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_334
timestamp 1644511149
transform 1 0 31832 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_342
timestamp 1644511149
transform 1 0 32568 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_347
timestamp 1644511149
transform 1 0 33028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_354
timestamp 1644511149
transform 1 0 33672 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1644511149
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_381
timestamp 1644511149
transform 1 0 36156 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_393
timestamp 1644511149
transform 1 0 37260 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_405
timestamp 1644511149
transform 1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_33
timestamp 1644511149
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_45
timestamp 1644511149
transform 1 0 5244 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1644511149
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_62
timestamp 1644511149
transform 1 0 6808 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_71
timestamp 1644511149
transform 1 0 7636 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_82
timestamp 1644511149
transform 1 0 8648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_91
timestamp 1644511149
transform 1 0 9476 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_97
timestamp 1644511149
transform 1 0 10028 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_103
timestamp 1644511149
transform 1 0 10580 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_116
timestamp 1644511149
transform 1 0 11776 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_120
timestamp 1644511149
transform 1 0 12144 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_126
timestamp 1644511149
transform 1 0 12696 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_133
timestamp 1644511149
transform 1 0 13340 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_143
timestamp 1644511149
transform 1 0 14260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1644511149
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_173
timestamp 1644511149
transform 1 0 17020 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_187
timestamp 1644511149
transform 1 0 18308 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_211
timestamp 1644511149
transform 1 0 20516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_229
timestamp 1644511149
transform 1 0 22172 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_235
timestamp 1644511149
transform 1 0 22724 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_252
timestamp 1644511149
transform 1 0 24288 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_256
timestamp 1644511149
transform 1 0 24656 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_299
timestamp 1644511149
transform 1 0 28612 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_307
timestamp 1644511149
transform 1 0 29348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_314
timestamp 1644511149
transform 1 0 29992 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_326
timestamp 1644511149
transform 1 0 31096 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 1644511149
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_342
timestamp 1644511149
transform 1 0 32568 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_356
timestamp 1644511149
transform 1 0 33856 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_362
timestamp 1644511149
transform 1 0 34408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_379
timestamp 1644511149
transform 1 0 35972 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1644511149
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1644511149
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_45
timestamp 1644511149
transform 1 0 5244 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_69
timestamp 1644511149
transform 1 0 7452 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_78
timestamp 1644511149
transform 1 0 8280 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_88
timestamp 1644511149
transform 1 0 9200 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_111
timestamp 1644511149
transform 1 0 11316 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1644511149
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_149
timestamp 1644511149
transform 1 0 14812 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_167
timestamp 1644511149
transform 1 0 16468 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_188
timestamp 1644511149
transform 1 0 18400 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_201
timestamp 1644511149
transform 1 0 19596 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_208
timestamp 1644511149
transform 1 0 20240 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_220
timestamp 1644511149
transform 1 0 21344 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_229
timestamp 1644511149
transform 1 0 22172 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_237
timestamp 1644511149
transform 1 0 22908 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_244
timestamp 1644511149
transform 1 0 23552 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_284
timestamp 1644511149
transform 1 0 27232 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_296
timestamp 1644511149
transform 1 0 28336 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1644511149
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_325
timestamp 1644511149
transform 1 0 31004 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_332
timestamp 1644511149
transform 1 0 31648 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_336
timestamp 1644511149
transform 1 0 32016 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_342
timestamp 1644511149
transform 1 0 32568 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_351
timestamp 1644511149
transform 1 0 33396 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_358
timestamp 1644511149
transform 1 0 34040 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_381
timestamp 1644511149
transform 1 0 36156 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_393
timestamp 1644511149
transform 1 0 37260 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_405
timestamp 1644511149
transform 1 0 38364 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_33
timestamp 1644511149
transform 1 0 4140 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_43
timestamp 1644511149
transform 1 0 5060 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1644511149
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_62
timestamp 1644511149
transform 1 0 6808 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_71
timestamp 1644511149
transform 1 0 7636 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_78
timestamp 1644511149
transform 1 0 8280 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_85
timestamp 1644511149
transform 1 0 8924 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_92
timestamp 1644511149
transform 1 0 9568 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_99
timestamp 1644511149
transform 1 0 10212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_134
timestamp 1644511149
transform 1 0 13432 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_146
timestamp 1644511149
transform 1 0 14536 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_152
timestamp 1644511149
transform 1 0 15088 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_162
timestamp 1644511149
transform 1 0 16008 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_190
timestamp 1644511149
transform 1 0 18584 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_212
timestamp 1644511149
transform 1 0 20608 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_241
timestamp 1644511149
transform 1 0 23276 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_250
timestamp 1644511149
transform 1 0 24104 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_257
timestamp 1644511149
transform 1 0 24748 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_263
timestamp 1644511149
transform 1 0 25300 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_269
timestamp 1644511149
transform 1 0 25852 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_277
timestamp 1644511149
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_302
timestamp 1644511149
transform 1 0 28888 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_310
timestamp 1644511149
transform 1 0 29624 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_326
timestamp 1644511149
transform 1 0 31096 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1644511149
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_359
timestamp 1644511149
transform 1 0 34132 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_379
timestamp 1644511149
transform 1 0 35972 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_386
timestamp 1644511149
transform 1 0 36616 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1644511149
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1644511149
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_45
timestamp 1644511149
transform 1 0 5244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_74
timestamp 1644511149
transform 1 0 7912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1644511149
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_88
timestamp 1644511149
transform 1 0 9200 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_110
timestamp 1644511149
transform 1 0 11224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_119
timestamp 1644511149
transform 1 0 12052 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_125
timestamp 1644511149
transform 1 0 12604 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_134
timestamp 1644511149
transform 1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_152
timestamp 1644511149
transform 1 0 15088 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_159
timestamp 1644511149
transform 1 0 15732 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_171
timestamp 1644511149
transform 1 0 16836 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_179
timestamp 1644511149
transform 1 0 17572 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_183
timestamp 1644511149
transform 1 0 17940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_205
timestamp 1644511149
transform 1 0 19964 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_211
timestamp 1644511149
transform 1 0 20516 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_220
timestamp 1644511149
transform 1 0 21344 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_231
timestamp 1644511149
transform 1 0 22356 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_239
timestamp 1644511149
transform 1 0 23092 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_244
timestamp 1644511149
transform 1 0 23552 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_261
timestamp 1644511149
transform 1 0 25116 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_269
timestamp 1644511149
transform 1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_275
timestamp 1644511149
transform 1 0 26404 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_287
timestamp 1644511149
transform 1 0 27508 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_291
timestamp 1644511149
transform 1 0 27876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_303
timestamp 1644511149
transform 1 0 28980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_313
timestamp 1644511149
transform 1 0 29900 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_322
timestamp 1644511149
transform 1 0 30728 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_331
timestamp 1644511149
transform 1 0 31556 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_340
timestamp 1644511149
transform 1 0 32384 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_360
timestamp 1644511149
transform 1 0 34224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_381
timestamp 1644511149
transform 1 0 36156 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_33
timestamp 1644511149
transform 1 0 4140 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_43
timestamp 1644511149
transform 1 0 5060 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1644511149
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_62
timestamp 1644511149
transform 1 0 6808 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_73
timestamp 1644511149
transform 1 0 7820 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_90
timestamp 1644511149
transform 1 0 9384 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_98
timestamp 1644511149
transform 1 0 10120 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1644511149
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1644511149
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_136
timestamp 1644511149
transform 1 0 13616 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_142
timestamp 1644511149
transform 1 0 14168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_159
timestamp 1644511149
transform 1 0 15732 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_186
timestamp 1644511149
transform 1 0 18216 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_193
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_206
timestamp 1644511149
transform 1 0 20056 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_215
timestamp 1644511149
transform 1 0 20884 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_229
timestamp 1644511149
transform 1 0 22172 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_236
timestamp 1644511149
transform 1 0 22816 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_245
timestamp 1644511149
transform 1 0 23644 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_253
timestamp 1644511149
transform 1 0 24380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_259
timestamp 1644511149
transform 1 0 24932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1644511149
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_288
timestamp 1644511149
transform 1 0 27600 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_296
timestamp 1644511149
transform 1 0 28336 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_303
timestamp 1644511149
transform 1 0 28980 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_315
timestamp 1644511149
transform 1 0 30084 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_323
timestamp 1644511149
transform 1 0 30820 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_332
timestamp 1644511149
transform 1 0 31648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_359
timestamp 1644511149
transform 1 0 34132 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_379
timestamp 1644511149
transform 1 0 35972 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_386
timestamp 1644511149
transform 1 0 36616 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_7
timestamp 1644511149
transform 1 0 1748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1644511149
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_45
timestamp 1644511149
transform 1 0 5244 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_60
timestamp 1644511149
transform 1 0 6624 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_69
timestamp 1644511149
transform 1 0 7452 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1644511149
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_90
timestamp 1644511149
transform 1 0 9384 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_102
timestamp 1644511149
transform 1 0 10488 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_113
timestamp 1644511149
transform 1 0 11500 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_125
timestamp 1644511149
transform 1 0 12604 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1644511149
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_155
timestamp 1644511149
transform 1 0 15364 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1644511149
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_167
timestamp 1644511149
transform 1 0 16468 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_176
timestamp 1644511149
transform 1 0 17296 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_187
timestamp 1644511149
transform 1 0 18308 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_213
timestamp 1644511149
transform 1 0 20700 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_228
timestamp 1644511149
transform 1 0 22080 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1644511149
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_259
timestamp 1644511149
transform 1 0 24932 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_267
timestamp 1644511149
transform 1 0 25668 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_272
timestamp 1644511149
transform 1 0 26128 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_300
timestamp 1644511149
transform 1 0 28704 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_314
timestamp 1644511149
transform 1 0 29992 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_324
timestamp 1644511149
transform 1 0 30912 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_342
timestamp 1644511149
transform 1 0 32568 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_351
timestamp 1644511149
transform 1 0 33396 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_358
timestamp 1644511149
transform 1 0 34040 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_33
timestamp 1644511149
transform 1 0 4140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_45
timestamp 1644511149
transform 1 0 5244 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1644511149
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_62
timestamp 1644511149
transform 1 0 6808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_76
timestamp 1644511149
transform 1 0 8096 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_83
timestamp 1644511149
transform 1 0 8740 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_95
timestamp 1644511149
transform 1 0 9844 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp 1644511149
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_118
timestamp 1644511149
transform 1 0 11960 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_126
timestamp 1644511149
transform 1 0 12696 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_136
timestamp 1644511149
transform 1 0 13616 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_145
timestamp 1644511149
transform 1 0 14444 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_157
timestamp 1644511149
transform 1 0 15548 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1644511149
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_173
timestamp 1644511149
transform 1 0 17020 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_177
timestamp 1644511149
transform 1 0 17388 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_195
timestamp 1644511149
transform 1 0 19044 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_207
timestamp 1644511149
transform 1 0 20148 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_219
timestamp 1644511149
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_234
timestamp 1644511149
transform 1 0 22632 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_240
timestamp 1644511149
transform 1 0 23184 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_251
timestamp 1644511149
transform 1 0 24196 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_260
timestamp 1644511149
transform 1 0 25024 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_266
timestamp 1644511149
transform 1 0 25576 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_284
timestamp 1644511149
transform 1 0 27232 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_290
timestamp 1644511149
transform 1 0 27784 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_307
timestamp 1644511149
transform 1 0 29348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_327
timestamp 1644511149
transform 1 0 31188 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_342
timestamp 1644511149
transform 1 0 32568 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_356
timestamp 1644511149
transform 1 0 33856 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_364
timestamp 1644511149
transform 1 0 34592 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_381
timestamp 1644511149
transform 1 0 36156 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1644511149
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_59
timestamp 1644511149
transform 1 0 6532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_66
timestamp 1644511149
transform 1 0 7176 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_78
timestamp 1644511149
transform 1 0 8280 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_93
timestamp 1644511149
transform 1 0 9660 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_101
timestamp 1644511149
transform 1 0 10396 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_112
timestamp 1644511149
transform 1 0 11408 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_124
timestamp 1644511149
transform 1 0 12512 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_149
timestamp 1644511149
transform 1 0 14812 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_154
timestamp 1644511149
transform 1 0 15272 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_162
timestamp 1644511149
transform 1 0 16008 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_170
timestamp 1644511149
transform 1 0 16744 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1644511149
transform 1 0 17480 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_190
timestamp 1644511149
transform 1 0 18584 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_202
timestamp 1644511149
transform 1 0 19688 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_214
timestamp 1644511149
transform 1 0 20792 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_234
timestamp 1644511149
transform 1 0 22632 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_243
timestamp 1644511149
transform 1 0 23460 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_257
timestamp 1644511149
transform 1 0 24748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_274
timestamp 1644511149
transform 1 0 26312 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_286
timestamp 1644511149
transform 1 0 27416 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_294
timestamp 1644511149
transform 1 0 28152 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_300
timestamp 1644511149
transform 1 0 28704 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_315
timestamp 1644511149
transform 1 0 30084 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_324
timestamp 1644511149
transform 1 0 30912 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_330
timestamp 1644511149
transform 1 0 31464 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_341
timestamp 1644511149
transform 1 0 32476 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_352
timestamp 1644511149
transform 1 0 33488 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_381
timestamp 1644511149
transform 1 0 36156 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_393
timestamp 1644511149
transform 1 0 37260 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_405
timestamp 1644511149
transform 1 0 38364 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1644511149
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1644511149
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1644511149
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_76
timestamp 1644511149
transform 1 0 8096 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_88
timestamp 1644511149
transform 1 0 9200 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1644511149
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_120
timestamp 1644511149
transform 1 0 12144 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_128
timestamp 1644511149
transform 1 0 12880 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_140
timestamp 1644511149
transform 1 0 13984 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_152
timestamp 1644511149
transform 1 0 15088 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_160
timestamp 1644511149
transform 1 0 15824 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_175
timestamp 1644511149
transform 1 0 17204 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1644511149
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_184
timestamp 1644511149
transform 1 0 18032 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_201
timestamp 1644511149
transform 1 0 19596 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_212
timestamp 1644511149
transform 1 0 20608 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1644511149
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_230
timestamp 1644511149
transform 1 0 22264 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_242
timestamp 1644511149
transform 1 0 23368 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_255
timestamp 1644511149
transform 1 0 24564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_259
timestamp 1644511149
transform 1 0 24932 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_264
timestamp 1644511149
transform 1 0 25392 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1644511149
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_305
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_317
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_325
timestamp 1644511149
transform 1 0 31004 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_333
timestamp 1644511149
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_342
timestamp 1644511149
transform 1 0 32568 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_346
timestamp 1644511149
transform 1 0 32936 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_357
timestamp 1644511149
transform 1 0 33948 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_369
timestamp 1644511149
transform 1 0 35052 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_381
timestamp 1644511149
transform 1 0 36156 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_389
timestamp 1644511149
transform 1 0 36892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_403
timestamp 1644511149
transform 1 0 38180 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_57
timestamp 1644511149
transform 1 0 6348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_63
timestamp 1644511149
transform 1 0 6900 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_75
timestamp 1644511149
transform 1 0 8004 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_79
timestamp 1644511149
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_108
timestamp 1644511149
transform 1 0 11040 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_120
timestamp 1644511149
transform 1 0 12144 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1644511149
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_151
timestamp 1644511149
transform 1 0 14996 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_155
timestamp 1644511149
transform 1 0 15364 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_164
timestamp 1644511149
transform 1 0 16192 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_176
timestamp 1644511149
transform 1 0 17296 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1644511149
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_213
timestamp 1644511149
transform 1 0 20700 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_225
timestamp 1644511149
transform 1 0 21804 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_234
timestamp 1644511149
transform 1 0 22632 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_242
timestamp 1644511149
transform 1 0 23368 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1644511149
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_261
timestamp 1644511149
transform 1 0 25116 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_273
timestamp 1644511149
transform 1 0 26220 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_284
timestamp 1644511149
transform 1 0 27232 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_293
timestamp 1644511149
transform 1 0 28060 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_305
timestamp 1644511149
transform 1 0 29164 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_337
timestamp 1644511149
transform 1 0 32108 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_341
timestamp 1644511149
transform 1 0 32476 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_347
timestamp 1644511149
transform 1 0 33028 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_353
timestamp 1644511149
transform 1 0 33580 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_359
timestamp 1644511149
transform 1 0 34132 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_375
timestamp 1644511149
transform 1 0 35604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_387
timestamp 1644511149
transform 1 0 36708 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_399
timestamp 1644511149
transform 1 0 37812 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_35
timestamp 1644511149
transform 1 0 4324 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_43
timestamp 1644511149
transform 1 0 5060 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1644511149
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_73
timestamp 1644511149
transform 1 0 7820 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_97
timestamp 1644511149
transform 1 0 10028 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1644511149
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_157
timestamp 1644511149
transform 1 0 15548 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1644511149
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_172
timestamp 1644511149
transform 1 0 16928 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_192
timestamp 1644511149
transform 1 0 18768 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_216
timestamp 1644511149
transform 1 0 20976 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_229
timestamp 1644511149
transform 1 0 22172 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_246
timestamp 1644511149
transform 1 0 23736 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_266
timestamp 1644511149
transform 1 0 25576 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1644511149
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_297
timestamp 1644511149
transform 1 0 28428 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_317
timestamp 1644511149
transform 1 0 30268 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_321
timestamp 1644511149
transform 1 0 30636 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_325
timestamp 1644511149
transform 1 0 31004 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_333
timestamp 1644511149
transform 1 0 31740 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_341
timestamp 1644511149
transform 1 0 32476 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_345
timestamp 1644511149
transform 1 0 32844 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_351
timestamp 1644511149
transform 1 0 33396 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_371
timestamp 1644511149
transform 1 0 35236 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_383
timestamp 1644511149
transform 1 0 36340 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_403
timestamp 1644511149
transform 1 0 38180 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_45
timestamp 1644511149
transform 1 0 5244 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_57
timestamp 1644511149
transform 1 0 6348 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_64
timestamp 1644511149
transform 1 0 6992 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_73
timestamp 1644511149
transform 1 0 7820 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1644511149
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_101
timestamp 1644511149
transform 1 0 10396 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_123
timestamp 1644511149
transform 1 0 12420 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_135
timestamp 1644511149
transform 1 0 13524 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_146
timestamp 1644511149
transform 1 0 14536 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_152
timestamp 1644511149
transform 1 0 15088 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_161
timestamp 1644511149
transform 1 0 15916 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_174
timestamp 1644511149
transform 1 0 17112 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_182
timestamp 1644511149
transform 1 0 17848 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1644511149
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_203
timestamp 1644511149
transform 1 0 19780 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_220
timestamp 1644511149
transform 1 0 21344 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_234
timestamp 1644511149
transform 1 0 22632 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_246
timestamp 1644511149
transform 1 0 23736 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_261
timestamp 1644511149
transform 1 0 25116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_273
timestamp 1644511149
transform 1 0 26220 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_282
timestamp 1644511149
transform 1 0 27048 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_294
timestamp 1644511149
transform 1 0 28152 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1644511149
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_335
timestamp 1644511149
transform 1 0 31924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_355
timestamp 1644511149
transform 1 0 33764 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_370
timestamp 1644511149
transform 1 0 35144 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_382
timestamp 1644511149
transform 1 0 36248 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_394
timestamp 1644511149
transform 1 0 37352 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_406
timestamp 1644511149
transform 1 0 38456 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_22
timestamp 1644511149
transform 1 0 3128 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_42
timestamp 1644511149
transform 1 0 4968 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_62
timestamp 1644511149
transform 1 0 6808 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_73
timestamp 1644511149
transform 1 0 7820 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_97
timestamp 1644511149
transform 1 0 10028 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_104
timestamp 1644511149
transform 1 0 10672 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_117
timestamp 1644511149
transform 1 0 11868 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_129
timestamp 1644511149
transform 1 0 12972 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_136
timestamp 1644511149
transform 1 0 13616 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_144
timestamp 1644511149
transform 1 0 14352 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_155
timestamp 1644511149
transform 1 0 15364 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1644511149
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_174
timestamp 1644511149
transform 1 0 17112 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_187
timestamp 1644511149
transform 1 0 18308 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_196
timestamp 1644511149
transform 1 0 19136 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_202
timestamp 1644511149
transform 1 0 19688 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_211
timestamp 1644511149
transform 1 0 20516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_233
timestamp 1644511149
transform 1 0 22540 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_239
timestamp 1644511149
transform 1 0 23092 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_251
timestamp 1644511149
transform 1 0 24196 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_257
timestamp 1644511149
transform 1 0 24748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_269
timestamp 1644511149
transform 1 0 25852 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 1644511149
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_286
timestamp 1644511149
transform 1 0 27416 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_325
timestamp 1644511149
transform 1 0 31004 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_333
timestamp 1644511149
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_345
timestamp 1644511149
transform 1 0 32844 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_353
timestamp 1644511149
transform 1 0 33580 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_368
timestamp 1644511149
transform 1 0 34960 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_380
timestamp 1644511149
transform 1 0 36064 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_45
timestamp 1644511149
transform 1 0 5244 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_59
timestamp 1644511149
transform 1 0 6532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_67
timestamp 1644511149
transform 1 0 7268 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_73
timestamp 1644511149
transform 1 0 7820 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1644511149
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_101
timestamp 1644511149
transform 1 0 10396 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_114
timestamp 1644511149
transform 1 0 11592 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_122
timestamp 1644511149
transform 1 0 12328 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_129
timestamp 1644511149
transform 1 0 12972 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_137
timestamp 1644511149
transform 1 0 13708 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_157
timestamp 1644511149
transform 1 0 15548 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_163
timestamp 1644511149
transform 1 0 16100 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_171
timestamp 1644511149
transform 1 0 16836 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_179
timestamp 1644511149
transform 1 0 17572 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1644511149
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_207
timestamp 1644511149
transform 1 0 20148 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_215
timestamp 1644511149
transform 1 0 20884 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_226
timestamp 1644511149
transform 1 0 21896 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_235
timestamp 1644511149
transform 1 0 22724 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_244
timestamp 1644511149
transform 1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_261
timestamp 1644511149
transform 1 0 25116 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_269
timestamp 1644511149
transform 1 0 25852 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_277
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_285
timestamp 1644511149
transform 1 0 27324 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_295
timestamp 1644511149
transform 1 0 28244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_314
timestamp 1644511149
transform 1 0 29992 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_336
timestamp 1644511149
transform 1 0 32016 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_348
timestamp 1644511149
transform 1 0 33120 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_352
timestamp 1644511149
transform 1 0 33488 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_358
timestamp 1644511149
transform 1 0 34040 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_33
timestamp 1644511149
transform 1 0 4140 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_37
timestamp 1644511149
transform 1 0 4508 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_44
timestamp 1644511149
transform 1 0 5152 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_67
timestamp 1644511149
transform 1 0 7268 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_76
timestamp 1644511149
transform 1 0 8096 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_83
timestamp 1644511149
transform 1 0 8740 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_87
timestamp 1644511149
transform 1 0 9108 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1644511149
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_129
timestamp 1644511149
transform 1 0 12972 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_141
timestamp 1644511149
transform 1 0 14076 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_147
timestamp 1644511149
transform 1 0 14628 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_153
timestamp 1644511149
transform 1 0 15180 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1644511149
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_173
timestamp 1644511149
transform 1 0 17020 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_209
timestamp 1644511149
transform 1 0 20332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_221
timestamp 1644511149
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_231
timestamp 1644511149
transform 1 0 22356 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_235
timestamp 1644511149
transform 1 0 22724 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_244
timestamp 1644511149
transform 1 0 23552 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_248
timestamp 1644511149
transform 1 0 23920 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_269
timestamp 1644511149
transform 1 0 25852 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_277
timestamp 1644511149
transform 1 0 26588 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_287
timestamp 1644511149
transform 1 0 27508 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_299
timestamp 1644511149
transform 1 0 28612 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_308
timestamp 1644511149
transform 1 0 29440 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_320
timestamp 1644511149
transform 1 0 30544 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_327
timestamp 1644511149
transform 1 0 31188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_344
timestamp 1644511149
transform 1 0 32752 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_352
timestamp 1644511149
transform 1 0 33488 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_369
timestamp 1644511149
transform 1 0 35052 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_381
timestamp 1644511149
transform 1 0 36156 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_389
timestamp 1644511149
transform 1 0 36892 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_79
timestamp 1644511149
transform 1 0 8372 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_130
timestamp 1644511149
transform 1 0 13064 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1644511149
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_163
timestamp 1644511149
transform 1 0 16100 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_183
timestamp 1644511149
transform 1 0 17940 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1644511149
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_220
timestamp 1644511149
transform 1 0 21344 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_228
timestamp 1644511149
transform 1 0 22080 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_248
timestamp 1644511149
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_263
timestamp 1644511149
transform 1 0 25300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_275
timestamp 1644511149
transform 1 0 26404 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_283
timestamp 1644511149
transform 1 0 27140 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_302
timestamp 1644511149
transform 1 0 28888 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_320
timestamp 1644511149
transform 1 0 30544 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_332
timestamp 1644511149
transform 1 0 31648 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_340
timestamp 1644511149
transform 1 0 32384 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_347
timestamp 1644511149
transform 1 0 33028 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_353
timestamp 1644511149
transform 1 0 33580 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1644511149
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_35
timestamp 1644511149
transform 1 0 4324 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_42
timestamp 1644511149
transform 1 0 4968 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1644511149
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_64
timestamp 1644511149
transform 1 0 6992 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_71
timestamp 1644511149
transform 1 0 7636 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_77
timestamp 1644511149
transform 1 0 8188 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_88
timestamp 1644511149
transform 1 0 9200 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_96
timestamp 1644511149
transform 1 0 9936 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_100
timestamp 1644511149
transform 1 0 10304 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_118
timestamp 1644511149
transform 1 0 11960 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_145
timestamp 1644511149
transform 1 0 14444 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_157
timestamp 1644511149
transform 1 0 15548 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_165
timestamp 1644511149
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_190
timestamp 1644511149
transform 1 0 18584 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_198
timestamp 1644511149
transform 1 0 19320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_219
timestamp 1644511149
transform 1 0 21252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_241
timestamp 1644511149
transform 1 0 23276 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_248
timestamp 1644511149
transform 1 0 23920 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_276
timestamp 1644511149
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_285
timestamp 1644511149
transform 1 0 27324 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_294
timestamp 1644511149
transform 1 0 28152 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_306
timestamp 1644511149
transform 1 0 29256 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_314
timestamp 1644511149
transform 1 0 29992 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1644511149
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_353
timestamp 1644511149
transform 1 0 33580 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_360
timestamp 1644511149
transform 1 0 34224 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_372
timestamp 1644511149
transform 1 0 35328 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_384
timestamp 1644511149
transform 1 0 36432 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_45
timestamp 1644511149
transform 1 0 5244 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_57
timestamp 1644511149
transform 1 0 6348 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_64
timestamp 1644511149
transform 1 0 6992 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_76
timestamp 1644511149
transform 1 0 8096 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1644511149
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_105
timestamp 1644511149
transform 1 0 10764 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_113
timestamp 1644511149
transform 1 0 11500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_125
timestamp 1644511149
transform 1 0 12604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_137
timestamp 1644511149
transform 1 0 13708 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_148
timestamp 1644511149
transform 1 0 14720 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_160
timestamp 1644511149
transform 1 0 15824 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_166
timestamp 1644511149
transform 1 0 16376 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_172
timestamp 1644511149
transform 1 0 16928 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_181
timestamp 1644511149
transform 1 0 17756 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_187
timestamp 1644511149
transform 1 0 18308 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1644511149
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_201
timestamp 1644511149
transform 1 0 19596 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_207
timestamp 1644511149
transform 1 0 20148 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_211
timestamp 1644511149
transform 1 0 20516 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_218
timestamp 1644511149
transform 1 0 21160 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_224
timestamp 1644511149
transform 1 0 21712 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_233
timestamp 1644511149
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1644511149
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_261
timestamp 1644511149
transform 1 0 25116 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_267
timestamp 1644511149
transform 1 0 25668 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_275
timestamp 1644511149
transform 1 0 26404 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_287
timestamp 1644511149
transform 1 0 27508 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_298
timestamp 1644511149
transform 1 0 28520 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_306
timestamp 1644511149
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_344
timestamp 1644511149
transform 1 0 32752 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_356
timestamp 1644511149
transform 1 0 33856 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_38
timestamp 1644511149
transform 1 0 4600 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_49
timestamp 1644511149
transform 1 0 5612 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_73
timestamp 1644511149
transform 1 0 7820 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_106
timestamp 1644511149
transform 1 0 10856 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_120
timestamp 1644511149
transform 1 0 12144 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_128
timestamp 1644511149
transform 1 0 12880 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_157
timestamp 1644511149
transform 1 0 15548 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_165
timestamp 1644511149
transform 1 0 16284 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_173
timestamp 1644511149
transform 1 0 17020 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_213
timestamp 1644511149
transform 1 0 20700 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 1644511149
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_235
timestamp 1644511149
transform 1 0 22724 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_243
timestamp 1644511149
transform 1 0 23460 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_255
timestamp 1644511149
transform 1 0 24564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_259
timestamp 1644511149
transform 1 0 24932 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_268
timestamp 1644511149
transform 1 0 25760 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_275
timestamp 1644511149
transform 1 0 26404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_303
timestamp 1644511149
transform 1 0 28980 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_307
timestamp 1644511149
transform 1 0 29348 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_313
timestamp 1644511149
transform 1 0 29900 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_326
timestamp 1644511149
transform 1 0 31096 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1644511149
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_46
timestamp 1644511149
transform 1 0 5336 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_54
timestamp 1644511149
transform 1 0 6072 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_71
timestamp 1644511149
transform 1 0 7636 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_80
timestamp 1644511149
transform 1 0 8464 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1644511149
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_98
timestamp 1644511149
transform 1 0 10120 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_106
timestamp 1644511149
transform 1 0 10856 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_114
timestamp 1644511149
transform 1 0 11592 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_127
timestamp 1644511149
transform 1 0 12788 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1644511149
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_177
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_185
timestamp 1644511149
transform 1 0 18124 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1644511149
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_205
timestamp 1644511149
transform 1 0 19964 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_213
timestamp 1644511149
transform 1 0 20700 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_225
timestamp 1644511149
transform 1 0 21804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_230
timestamp 1644511149
transform 1 0 22264 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_240
timestamp 1644511149
transform 1 0 23184 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1644511149
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_258
timestamp 1644511149
transform 1 0 24840 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_266
timestamp 1644511149
transform 1 0 25576 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_272
timestamp 1644511149
transform 1 0 26128 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_284
timestamp 1644511149
transform 1 0 27232 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_299
timestamp 1644511149
transform 1 0 28612 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_325
timestamp 1644511149
transform 1 0 31004 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_345
timestamp 1644511149
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_35
timestamp 1644511149
transform 1 0 4324 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_40
timestamp 1644511149
transform 1 0 4784 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1644511149
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_68
timestamp 1644511149
transform 1 0 7360 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_80
timestamp 1644511149
transform 1 0 8464 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_95
timestamp 1644511149
transform 1 0 9844 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_103
timestamp 1644511149
transform 1 0 10580 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_108
timestamp 1644511149
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_129
timestamp 1644511149
transform 1 0 12972 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_141
timestamp 1644511149
transform 1 0 14076 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1644511149
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_177
timestamp 1644511149
transform 1 0 17388 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_187
timestamp 1644511149
transform 1 0 18308 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_196
timestamp 1644511149
transform 1 0 19136 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_218
timestamp 1644511149
transform 1 0 21160 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_230
timestamp 1644511149
transform 1 0 22264 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_238
timestamp 1644511149
transform 1 0 23000 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_246
timestamp 1644511149
transform 1 0 23736 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_257
timestamp 1644511149
transform 1 0 24748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_265
timestamp 1644511149
transform 1 0 25484 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_269
timestamp 1644511149
transform 1 0 25852 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_275
timestamp 1644511149
transform 1 0 26404 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_297
timestamp 1644511149
transform 1 0 28428 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_313
timestamp 1644511149
transform 1 0 29900 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_323
timestamp 1644511149
transform 1 0 30820 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_330
timestamp 1644511149
transform 1 0 31464 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_50
timestamp 1644511149
transform 1 0 5704 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_58
timestamp 1644511149
transform 1 0 6440 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_64
timestamp 1644511149
transform 1 0 6992 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_76
timestamp 1644511149
transform 1 0 8096 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_89
timestamp 1644511149
transform 1 0 9292 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_100
timestamp 1644511149
transform 1 0 10304 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_115
timestamp 1644511149
transform 1 0 11684 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_125
timestamp 1644511149
transform 1 0 12604 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_130
timestamp 1644511149
transform 1 0 13064 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1644511149
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_163
timestamp 1644511149
transform 1 0 16100 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_167
timestamp 1644511149
transform 1 0 16468 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_173
timestamp 1644511149
transform 1 0 17020 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_185
timestamp 1644511149
transform 1 0 18124 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_193
timestamp 1644511149
transform 1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_217
timestamp 1644511149
transform 1 0 21068 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_222
timestamp 1644511149
transform 1 0 21528 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_230
timestamp 1644511149
transform 1 0 22264 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1644511149
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_269
timestamp 1644511149
transform 1 0 25852 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_281
timestamp 1644511149
transform 1 0 26956 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_298
timestamp 1644511149
transform 1 0 28520 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 1644511149
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_317
timestamp 1644511149
transform 1 0 30268 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_326
timestamp 1644511149
transform 1 0 31096 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_338
timestamp 1644511149
transform 1 0 32200 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_350
timestamp 1644511149
transform 1 0 33304 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 1644511149
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_47
timestamp 1644511149
transform 1 0 5428 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_62
timestamp 1644511149
transform 1 0 6808 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_70
timestamp 1644511149
transform 1 0 7544 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_77
timestamp 1644511149
transform 1 0 8188 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_101
timestamp 1644511149
transform 1 0 10396 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp 1644511149
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_147
timestamp 1644511149
transform 1 0 14628 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_155
timestamp 1644511149
transform 1 0 15364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_162
timestamp 1644511149
transform 1 0 16008 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_187
timestamp 1644511149
transform 1 0 18308 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_199
timestamp 1644511149
transform 1 0 19412 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_211
timestamp 1644511149
transform 1 0 20516 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_219
timestamp 1644511149
transform 1 0 21252 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_249
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_264
timestamp 1644511149
transform 1 0 25392 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1644511149
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_297
timestamp 1644511149
transform 1 0 28428 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_309
timestamp 1644511149
transform 1 0 29532 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_323
timestamp 1644511149
transform 1 0 30820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_57
timestamp 1644511149
transform 1 0 6348 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_63
timestamp 1644511149
transform 1 0 6900 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp 1644511149
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_101
timestamp 1644511149
transform 1 0 10396 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_126
timestamp 1644511149
transform 1 0 12696 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_136
timestamp 1644511149
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_158
timestamp 1644511149
transform 1 0 15640 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_170
timestamp 1644511149
transform 1 0 16744 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_182
timestamp 1644511149
transform 1 0 17848 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1644511149
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_207
timestamp 1644511149
transform 1 0 20148 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_211
timestamp 1644511149
transform 1 0 20516 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_228
timestamp 1644511149
transform 1 0 22080 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_242
timestamp 1644511149
transform 1 0 23368 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1644511149
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_302
timestamp 1644511149
transform 1 0 28888 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_313
timestamp 1644511149
transform 1 0 29900 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_330
timestamp 1644511149
transform 1 0 31464 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_342
timestamp 1644511149
transform 1 0 32568 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_354
timestamp 1644511149
transform 1 0 33672 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_362
timestamp 1644511149
transform 1 0 34408 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_35
timestamp 1644511149
transform 1 0 4324 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_52
timestamp 1644511149
transform 1 0 5888 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_62
timestamp 1644511149
transform 1 0 6808 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_76
timestamp 1644511149
transform 1 0 8096 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_83
timestamp 1644511149
transform 1 0 8740 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_91
timestamp 1644511149
transform 1 0 9476 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_97
timestamp 1644511149
transform 1 0 10028 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_104
timestamp 1644511149
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_133
timestamp 1644511149
transform 1 0 13340 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_143
timestamp 1644511149
transform 1 0 14260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_163
timestamp 1644511149
transform 1 0 16100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_177
timestamp 1644511149
transform 1 0 17388 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_186
timestamp 1644511149
transform 1 0 18216 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_206
timestamp 1644511149
transform 1 0 20056 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1644511149
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_233
timestamp 1644511149
transform 1 0 22540 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_239
timestamp 1644511149
transform 1 0 23092 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_245
timestamp 1644511149
transform 1 0 23644 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_252
timestamp 1644511149
transform 1 0 24288 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_259
timestamp 1644511149
transform 1 0 24932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_263
timestamp 1644511149
transform 1 0 25300 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_272
timestamp 1644511149
transform 1 0 26128 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_285
timestamp 1644511149
transform 1 0 27324 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_294
timestamp 1644511149
transform 1 0 28152 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_306
timestamp 1644511149
transform 1 0 29256 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_45_328
timestamp 1644511149
transform 1 0 31280 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_45
timestamp 1644511149
transform 1 0 5244 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_62
timestamp 1644511149
transform 1 0 6808 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_70
timestamp 1644511149
transform 1 0 7544 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_101
timestamp 1644511149
transform 1 0 10396 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_106
timestamp 1644511149
transform 1 0 10856 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_118
timestamp 1644511149
transform 1 0 11960 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_122
timestamp 1644511149
transform 1 0 12328 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_128
timestamp 1644511149
transform 1 0 12880 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1644511149
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_145
timestamp 1644511149
transform 1 0 14444 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_151
timestamp 1644511149
transform 1 0 14996 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_171
timestamp 1644511149
transform 1 0 16836 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_181
timestamp 1644511149
transform 1 0 17756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_193
timestamp 1644511149
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_205
timestamp 1644511149
transform 1 0 19964 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_218
timestamp 1644511149
transform 1 0 21160 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_230
timestamp 1644511149
transform 1 0 22264 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_240
timestamp 1644511149
transform 1 0 23184 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1644511149
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_259
timestamp 1644511149
transform 1 0 24932 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_267
timestamp 1644511149
transform 1 0 25668 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_276
timestamp 1644511149
transform 1 0 26496 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_285
timestamp 1644511149
transform 1 0 27324 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_298
timestamp 1644511149
transform 1 0 28520 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_306
timestamp 1644511149
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_317
timestamp 1644511149
transform 1 0 30268 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_329
timestamp 1644511149
transform 1 0 31372 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_341
timestamp 1644511149
transform 1 0 32476 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_353
timestamp 1644511149
transform 1 0 33580 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_361
timestamp 1644511149
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_63
timestamp 1644511149
transform 1 0 6900 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_83
timestamp 1644511149
transform 1 0 8740 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_103
timestamp 1644511149
transform 1 0 10580 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_130
timestamp 1644511149
transform 1 0 13064 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_138
timestamp 1644511149
transform 1 0 13800 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_146
timestamp 1644511149
transform 1 0 14536 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_152
timestamp 1644511149
transform 1 0 15088 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1644511149
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_187
timestamp 1644511149
transform 1 0 18308 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_197
timestamp 1644511149
transform 1 0 19228 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_205
timestamp 1644511149
transform 1 0 19964 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_213
timestamp 1644511149
transform 1 0 20700 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_219
timestamp 1644511149
transform 1 0 21252 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_242
timestamp 1644511149
transform 1 0 23368 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_246
timestamp 1644511149
transform 1 0 23736 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_254
timestamp 1644511149
transform 1 0 24472 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1644511149
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_326
timestamp 1644511149
transform 1 0 31096 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_334
timestamp 1644511149
transform 1 0 31832 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_361
timestamp 1644511149
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_373
timestamp 1644511149
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1644511149
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_47
timestamp 1644511149
transform 1 0 5428 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_68
timestamp 1644511149
transform 1 0 7360 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_101
timestamp 1644511149
transform 1 0 10396 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_122
timestamp 1644511149
transform 1 0 12328 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_134
timestamp 1644511149
transform 1 0 13432 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_145
timestamp 1644511149
transform 1 0 14444 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_154
timestamp 1644511149
transform 1 0 15272 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_158
timestamp 1644511149
transform 1 0 15640 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_175
timestamp 1644511149
transform 1 0 17204 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_183
timestamp 1644511149
transform 1 0 17940 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_191
timestamp 1644511149
transform 1 0 18676 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_201
timestamp 1644511149
transform 1 0 19596 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_242
timestamp 1644511149
transform 1 0 23368 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1644511149
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_258
timestamp 1644511149
transform 1 0 24840 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_262
timestamp 1644511149
transform 1 0 25208 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_268
timestamp 1644511149
transform 1 0 25760 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_284
timestamp 1644511149
transform 1 0 27232 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_294
timestamp 1644511149
transform 1 0 28152 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_302
timestamp 1644511149
transform 1 0 28888 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_319
timestamp 1644511149
transform 1 0 30452 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_325
timestamp 1644511149
transform 1 0 31004 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_346
timestamp 1644511149
transform 1 0 32936 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_358
timestamp 1644511149
transform 1 0 34040 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_35
timestamp 1644511149
transform 1 0 4324 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_52
timestamp 1644511149
transform 1 0 5888 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_62
timestamp 1644511149
transform 1 0 6808 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_70
timestamp 1644511149
transform 1 0 7544 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_82
timestamp 1644511149
transform 1 0 8648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_102
timestamp 1644511149
transform 1 0 10488 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1644511149
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_122
timestamp 1644511149
transform 1 0 12328 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_142
timestamp 1644511149
transform 1 0 14168 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_162
timestamp 1644511149
transform 1 0 16008 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_177
timestamp 1644511149
transform 1 0 17388 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_185
timestamp 1644511149
transform 1 0 18124 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_213
timestamp 1644511149
transform 1 0 20700 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_221
timestamp 1644511149
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_241
timestamp 1644511149
transform 1 0 23276 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_250
timestamp 1644511149
transform 1 0 24104 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_258
timestamp 1644511149
transform 1 0 24840 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_272
timestamp 1644511149
transform 1 0 26128 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_297
timestamp 1644511149
transform 1 0 28428 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_306
timestamp 1644511149
transform 1 0 29256 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_318
timestamp 1644511149
transform 1 0 30360 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_330
timestamp 1644511149
transform 1 0 31464 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_37
timestamp 1644511149
transform 1 0 4508 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_43
timestamp 1644511149
transform 1 0 5060 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_52
timestamp 1644511149
transform 1 0 5888 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_59
timestamp 1644511149
transform 1 0 6532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_71
timestamp 1644511149
transform 1 0 7636 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_75
timestamp 1644511149
transform 1 0 8004 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_94
timestamp 1644511149
transform 1 0 9752 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_114
timestamp 1644511149
transform 1 0 11592 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_123
timestamp 1644511149
transform 1 0 12420 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_132
timestamp 1644511149
transform 1 0 13248 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_146
timestamp 1644511149
transform 1 0 14536 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_158
timestamp 1644511149
transform 1 0 15640 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_170
timestamp 1644511149
transform 1 0 16744 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_182
timestamp 1644511149
transform 1 0 17848 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1644511149
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_202
timestamp 1644511149
transform 1 0 19688 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_210
timestamp 1644511149
transform 1 0 20424 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_232
timestamp 1644511149
transform 1 0 22448 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_238
timestamp 1644511149
transform 1 0 23000 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_247
timestamp 1644511149
transform 1 0 23828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_257
timestamp 1644511149
transform 1 0 24748 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_263
timestamp 1644511149
transform 1 0 25300 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_280
timestamp 1644511149
transform 1 0 26864 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_286
timestamp 1644511149
transform 1 0 27416 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_303
timestamp 1644511149
transform 1 0 28980 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_331
timestamp 1644511149
transform 1 0 31556 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_351
timestamp 1644511149
transform 1 0 33396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_77
timestamp 1644511149
transform 1 0 8188 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_89
timestamp 1644511149
transform 1 0 9292 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_101
timestamp 1644511149
transform 1 0 10396 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_109
timestamp 1644511149
transform 1 0 11132 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_154
timestamp 1644511149
transform 1 0 15272 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1644511149
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_177
timestamp 1644511149
transform 1 0 17388 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_187
timestamp 1644511149
transform 1 0 18308 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_194
timestamp 1644511149
transform 1 0 18952 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_206
timestamp 1644511149
transform 1 0 20056 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_213
timestamp 1644511149
transform 1 0 20700 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_221
timestamp 1644511149
transform 1 0 21436 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_231
timestamp 1644511149
transform 1 0 22356 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_236
timestamp 1644511149
transform 1 0 22816 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_257
timestamp 1644511149
transform 1 0 24748 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_289
timestamp 1644511149
transform 1 0 27692 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_297
timestamp 1644511149
transform 1 0 28428 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_309
timestamp 1644511149
transform 1 0 29532 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_321
timestamp 1644511149
transform 1 0 30636 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_333
timestamp 1644511149
transform 1 0 31740 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1644511149
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_58
timestamp 1644511149
transform 1 0 6440 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_64
timestamp 1644511149
transform 1 0 6992 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_68
timestamp 1644511149
transform 1 0 7360 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_117
timestamp 1644511149
transform 1 0 11868 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_127
timestamp 1644511149
transform 1 0 12788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_149
timestamp 1644511149
transform 1 0 14812 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_155
timestamp 1644511149
transform 1 0 15364 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_172
timestamp 1644511149
transform 1 0 16928 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1644511149
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_205
timestamp 1644511149
transform 1 0 19964 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_217
timestamp 1644511149
transform 1 0 21068 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_229
timestamp 1644511149
transform 1 0 22172 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_237
timestamp 1644511149
transform 1 0 22908 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1644511149
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_260
timestamp 1644511149
transform 1 0 25024 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_272
timestamp 1644511149
transform 1 0 26128 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_284
timestamp 1644511149
transform 1 0 27232 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_298
timestamp 1644511149
transform 1 0 28520 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_306
timestamp 1644511149
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_345
timestamp 1644511149
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1644511149
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_52
timestamp 1644511149
transform 1 0 5888 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_62
timestamp 1644511149
transform 1 0 6808 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_82
timestamp 1644511149
transform 1 0 8648 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_90
timestamp 1644511149
transform 1 0 9384 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_100
timestamp 1644511149
transform 1 0 10304 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_129
timestamp 1644511149
transform 1 0 12972 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_139
timestamp 1644511149
transform 1 0 13892 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_159
timestamp 1644511149
transform 1 0 15732 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_174
timestamp 1644511149
transform 1 0 17112 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_182
timestamp 1644511149
transform 1 0 17848 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_188
timestamp 1644511149
transform 1 0 18400 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_198
timestamp 1644511149
transform 1 0 19320 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_210
timestamp 1644511149
transform 1 0 20424 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1644511149
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_233
timestamp 1644511149
transform 1 0 22540 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_239
timestamp 1644511149
transform 1 0 23092 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_248
timestamp 1644511149
transform 1 0 23920 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_256
timestamp 1644511149
transform 1 0 24656 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_275
timestamp 1644511149
transform 1 0 26404 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_295
timestamp 1644511149
transform 1 0 28244 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_301
timestamp 1644511149
transform 1 0 28796 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_318
timestamp 1644511149
transform 1 0 30360 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_325
timestamp 1644511149
transform 1 0 31004 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_333
timestamp 1644511149
transform 1 0 31740 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_373
timestamp 1644511149
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_58
timestamp 1644511149
transform 1 0 6440 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_80
timestamp 1644511149
transform 1 0 8464 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_104
timestamp 1644511149
transform 1 0 10672 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_116
timestamp 1644511149
transform 1 0 11776 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_136
timestamp 1644511149
transform 1 0 13616 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_147
timestamp 1644511149
transform 1 0 14628 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_155
timestamp 1644511149
transform 1 0 15364 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_178
timestamp 1644511149
transform 1 0 17480 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_190
timestamp 1644511149
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_205
timestamp 1644511149
transform 1 0 19964 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_211
timestamp 1644511149
transform 1 0 20516 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_228
timestamp 1644511149
transform 1 0 22080 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp 1644511149
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_261
timestamp 1644511149
transform 1 0 25116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_272
timestamp 1644511149
transform 1 0 26128 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_284
timestamp 1644511149
transform 1 0 27232 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_294
timestamp 1644511149
transform 1 0 28152 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_306
timestamp 1644511149
transform 1 0 29256 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_322
timestamp 1644511149
transform 1 0 30728 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_329
timestamp 1644511149
transform 1 0 31372 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_341
timestamp 1644511149
transform 1 0 32476 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_353
timestamp 1644511149
transform 1 0 33580 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_361
timestamp 1644511149
transform 1 0 34316 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_47
timestamp 1644511149
transform 1 0 5428 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1644511149
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_60
timestamp 1644511149
transform 1 0 6624 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_75
timestamp 1644511149
transform 1 0 8004 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_87
timestamp 1644511149
transform 1 0 9108 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_91
timestamp 1644511149
transform 1 0 9476 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_108
timestamp 1644511149
transform 1 0 11040 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_118
timestamp 1644511149
transform 1 0 11960 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_126
timestamp 1644511149
transform 1 0 12696 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_145
timestamp 1644511149
transform 1 0 14444 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_156
timestamp 1644511149
transform 1 0 15456 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_164
timestamp 1644511149
transform 1 0 16192 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_179
timestamp 1644511149
transform 1 0 17572 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_187
timestamp 1644511149
transform 1 0 18308 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_204
timestamp 1644511149
transform 1 0 19872 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_212
timestamp 1644511149
transform 1 0 20608 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_233
timestamp 1644511149
transform 1 0 22540 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_245
timestamp 1644511149
transform 1 0 23644 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_55_256
timestamp 1644511149
transform 1 0 24656 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_262
timestamp 1644511149
transform 1 0 25208 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_269
timestamp 1644511149
transform 1 0 25852 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_277
timestamp 1644511149
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_290
timestamp 1644511149
transform 1 0 27784 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_300
timestamp 1644511149
transform 1 0 28704 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_312
timestamp 1644511149
transform 1 0 29808 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_332
timestamp 1644511149
transform 1 0 31648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_89
timestamp 1644511149
transform 1 0 9292 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_101
timestamp 1644511149
transform 1 0 10396 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_110
timestamp 1644511149
transform 1 0 11224 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_118
timestamp 1644511149
transform 1 0 11960 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_127
timestamp 1644511149
transform 1 0 12788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_157
timestamp 1644511149
transform 1 0 15548 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_163
timestamp 1644511149
transform 1 0 16100 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_174
timestamp 1644511149
transform 1 0 17112 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_178
timestamp 1644511149
transform 1 0 17480 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_203
timestamp 1644511149
transform 1 0 19780 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_211
timestamp 1644511149
transform 1 0 20516 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_223
timestamp 1644511149
transform 1 0 21620 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_232
timestamp 1644511149
transform 1 0 22448 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_240
timestamp 1644511149
transform 1 0 23184 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1644511149
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_275
timestamp 1644511149
transform 1 0 26404 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_287
timestamp 1644511149
transform 1 0 27508 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_304
timestamp 1644511149
transform 1 0 29072 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_317
timestamp 1644511149
transform 1 0 30268 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_323
timestamp 1644511149
transform 1 0 30820 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_335
timestamp 1644511149
transform 1 0 31924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_347
timestamp 1644511149
transform 1 0 33028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_359
timestamp 1644511149
transform 1 0 34132 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_102
timestamp 1644511149
transform 1 0 10488 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_110
timestamp 1644511149
transform 1 0 11224 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_117
timestamp 1644511149
transform 1 0 11868 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_126
timestamp 1644511149
transform 1 0 12696 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_134
timestamp 1644511149
transform 1 0 13432 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_144
timestamp 1644511149
transform 1 0 14352 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_156
timestamp 1644511149
transform 1 0 15456 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_163
timestamp 1644511149
transform 1 0 16100 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_179
timestamp 1644511149
transform 1 0 17572 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_207
timestamp 1644511149
transform 1 0 20148 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_219
timestamp 1644511149
transform 1 0 21252 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_245
timestamp 1644511149
transform 1 0 23644 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_253
timestamp 1644511149
transform 1 0 24380 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_259
timestamp 1644511149
transform 1 0 24932 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_276
timestamp 1644511149
transform 1 0 26496 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_303
timestamp 1644511149
transform 1 0 28980 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_311
timestamp 1644511149
transform 1 0 29716 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_315
timestamp 1644511149
transform 1 0 30084 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_319
timestamp 1644511149
transform 1 0 30452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_331
timestamp 1644511149
transform 1 0 31556 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_89
timestamp 1644511149
transform 1 0 9292 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_98
timestamp 1644511149
transform 1 0 10120 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_112
timestamp 1644511149
transform 1 0 11408 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_129
timestamp 1644511149
transform 1 0 12972 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_136
timestamp 1644511149
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_149
timestamp 1644511149
transform 1 0 14812 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_160
timestamp 1644511149
transform 1 0 15824 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_173
timestamp 1644511149
transform 1 0 17020 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_187
timestamp 1644511149
transform 1 0 18308 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_206
timestamp 1644511149
transform 1 0 20056 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_219
timestamp 1644511149
transform 1 0 21252 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_232
timestamp 1644511149
transform 1 0 22448 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_240
timestamp 1644511149
transform 1 0 23184 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1644511149
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_256
timestamp 1644511149
transform 1 0 24656 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_264
timestamp 1644511149
transform 1 0 25392 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_287
timestamp 1644511149
transform 1 0 27508 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_294
timestamp 1644511149
transform 1 0 28152 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_306
timestamp 1644511149
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_312
timestamp 1644511149
transform 1 0 29808 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_323
timestamp 1644511149
transform 1 0 30820 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_330
timestamp 1644511149
transform 1 0 31464 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_342
timestamp 1644511149
transform 1 0 32568 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_354
timestamp 1644511149
transform 1 0 33672 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_362
timestamp 1644511149
transform 1 0 34408 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_90
timestamp 1644511149
transform 1 0 9384 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_104
timestamp 1644511149
transform 1 0 10672 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_128
timestamp 1644511149
transform 1 0 12880 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_145
timestamp 1644511149
transform 1 0 14444 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_163
timestamp 1644511149
transform 1 0 16100 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_177
timestamp 1644511149
transform 1 0 17388 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_189
timestamp 1644511149
transform 1 0 18492 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_199
timestamp 1644511149
transform 1 0 19412 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_203
timestamp 1644511149
transform 1 0 19780 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_212
timestamp 1644511149
transform 1 0 20608 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_216
timestamp 1644511149
transform 1 0 20976 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_220
timestamp 1644511149
transform 1 0 21344 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_230
timestamp 1644511149
transform 1 0 22264 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_241
timestamp 1644511149
transform 1 0 23276 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_248
timestamp 1644511149
transform 1 0 23920 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_260
timestamp 1644511149
transform 1 0 25024 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_266
timestamp 1644511149
transform 1 0 25576 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_270
timestamp 1644511149
transform 1 0 25944 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_278
timestamp 1644511149
transform 1 0 26680 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_300
timestamp 1644511149
transform 1 0 28704 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_312
timestamp 1644511149
transform 1 0 29808 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_332
timestamp 1644511149
transform 1 0 31648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_93
timestamp 1644511149
transform 1 0 9660 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_103
timestamp 1644511149
transform 1 0 10580 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_112
timestamp 1644511149
transform 1 0 11408 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_119
timestamp 1644511149
transform 1 0 12052 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_127
timestamp 1644511149
transform 1 0 12788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_150
timestamp 1644511149
transform 1 0 14904 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_162
timestamp 1644511149
transform 1 0 16008 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_171
timestamp 1644511149
transform 1 0 16836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_186
timestamp 1644511149
transform 1 0 18216 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_194
timestamp 1644511149
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_200
timestamp 1644511149
transform 1 0 19504 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_212
timestamp 1644511149
transform 1 0 20608 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_216
timestamp 1644511149
transform 1 0 20976 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_226
timestamp 1644511149
transform 1 0 21896 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_241
timestamp 1644511149
transform 1 0 23276 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_248
timestamp 1644511149
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_259
timestamp 1644511149
transform 1 0 24932 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_266
timestamp 1644511149
transform 1 0 25576 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_273
timestamp 1644511149
transform 1 0 26220 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_285
timestamp 1644511149
transform 1 0 27324 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_297
timestamp 1644511149
transform 1 0 28428 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_304
timestamp 1644511149
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_319
timestamp 1644511149
transform 1 0 30452 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_328
timestamp 1644511149
transform 1 0 31280 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_340
timestamp 1644511149
transform 1 0 32384 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_352
timestamp 1644511149
transform 1 0 33488 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1644511149
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_100
timestamp 1644511149
transform 1 0 10304 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_129
timestamp 1644511149
transform 1 0 12972 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_185
timestamp 1644511149
transform 1 0 18124 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_198
timestamp 1644511149
transform 1 0 19320 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_207
timestamp 1644511149
transform 1 0 20148 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_214
timestamp 1644511149
transform 1 0 20792 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1644511149
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_233
timestamp 1644511149
transform 1 0 22540 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_61_255
timestamp 1644511149
transform 1 0 24564 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_263
timestamp 1644511149
transform 1 0 25300 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_272
timestamp 1644511149
transform 1 0 26128 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_289
timestamp 1644511149
transform 1 0 27692 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_296
timestamp 1644511149
transform 1 0 28336 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_303
timestamp 1644511149
transform 1 0 28980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_313
timestamp 1644511149
transform 1 0 29900 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_317
timestamp 1644511149
transform 1 0 30268 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_323
timestamp 1644511149
transform 1 0 30820 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_113
timestamp 1644511149
transform 1 0 11500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_117
timestamp 1644511149
transform 1 0 11868 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_129
timestamp 1644511149
transform 1 0 12972 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_134
timestamp 1644511149
transform 1 0 13432 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_161
timestamp 1644511149
transform 1 0 15916 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_166
timestamp 1644511149
transform 1 0 16376 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_174
timestamp 1644511149
transform 1 0 17112 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_62_187
timestamp 1644511149
transform 1 0 18308 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_204
timestamp 1644511149
transform 1 0 19872 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_212
timestamp 1644511149
transform 1 0 20608 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_227
timestamp 1644511149
transform 1 0 21988 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_233
timestamp 1644511149
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1644511149
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_270
timestamp 1644511149
transform 1 0 25944 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_277
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_289
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_62_300
timestamp 1644511149
transform 1 0 28704 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1644511149
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_89
timestamp 1644511149
transform 1 0 9292 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_108
timestamp 1644511149
transform 1 0 11040 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_118
timestamp 1644511149
transform 1 0 11960 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_136
timestamp 1644511149
transform 1 0 13616 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_143
timestamp 1644511149
transform 1 0 14260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_155
timestamp 1644511149
transform 1 0 15364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_164
timestamp 1644511149
transform 1 0 16192 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_174
timestamp 1644511149
transform 1 0 17112 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_192
timestamp 1644511149
transform 1 0 18768 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_201
timestamp 1644511149
transform 1 0 19596 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_214
timestamp 1644511149
transform 1 0 20792 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1644511149
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_232
timestamp 1644511149
transform 1 0 22448 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_241
timestamp 1644511149
transform 1 0 23276 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_248
timestamp 1644511149
transform 1 0 23920 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_255
timestamp 1644511149
transform 1 0 24564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_259
timestamp 1644511149
transform 1 0 24932 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1644511149
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_287
timestamp 1644511149
transform 1 0 27508 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_291
timestamp 1644511149
transform 1 0 27876 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_302
timestamp 1644511149
transform 1 0 28888 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_314
timestamp 1644511149
transform 1 0 29992 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_326
timestamp 1644511149
transform 1 0 31096 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_334
timestamp 1644511149
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_102
timestamp 1644511149
transform 1 0 10488 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_114
timestamp 1644511149
transform 1 0 11592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_122
timestamp 1644511149
transform 1 0 12328 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_128
timestamp 1644511149
transform 1 0 12880 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_135
timestamp 1644511149
transform 1 0 13524 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_157
timestamp 1644511149
transform 1 0 15548 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_169
timestamp 1644511149
transform 1 0 16652 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_187
timestamp 1644511149
transform 1 0 18308 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_222
timestamp 1644511149
transform 1 0 21528 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_234
timestamp 1644511149
transform 1 0 22632 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_240
timestamp 1644511149
transform 1 0 23184 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 1644511149
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_260
timestamp 1644511149
transform 1 0 25024 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_280
timestamp 1644511149
transform 1 0 26864 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_304
timestamp 1644511149
transform 1 0 29072 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_129
timestamp 1644511149
transform 1 0 12972 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_144
timestamp 1644511149
transform 1 0 14352 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_153
timestamp 1644511149
transform 1 0 15180 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_165
timestamp 1644511149
transform 1 0 16284 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_65_179
timestamp 1644511149
transform 1 0 17572 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_185
timestamp 1644511149
transform 1 0 18124 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_197
timestamp 1644511149
transform 1 0 19228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_201
timestamp 1644511149
transform 1 0 19596 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_208
timestamp 1644511149
transform 1 0 20240 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_220
timestamp 1644511149
transform 1 0 21344 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_230
timestamp 1644511149
transform 1 0 22264 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_242
timestamp 1644511149
transform 1 0 23368 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_254
timestamp 1644511149
transform 1 0 24472 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_260
timestamp 1644511149
transform 1 0 25024 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_264
timestamp 1644511149
transform 1 0 25392 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_276
timestamp 1644511149
transform 1 0 26496 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_291
timestamp 1644511149
transform 1 0 27876 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_301
timestamp 1644511149
transform 1 0 28796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_310
timestamp 1644511149
transform 1 0 29624 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_322
timestamp 1644511149
transform 1 0 30728 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_334
timestamp 1644511149
transform 1 0 31832 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_103
timestamp 1644511149
transform 1 0 10580 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_124
timestamp 1644511149
transform 1 0 12512 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_128
timestamp 1644511149
transform 1 0 12880 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_135
timestamp 1644511149
transform 1 0 13524 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_144
timestamp 1644511149
transform 1 0 14352 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_161
timestamp 1644511149
transform 1 0 15916 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_172
timestamp 1644511149
transform 1 0 16928 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_184
timestamp 1644511149
transform 1 0 18032 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_206
timestamp 1644511149
transform 1 0 20056 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_214
timestamp 1644511149
transform 1 0 20792 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_224
timestamp 1644511149
transform 1 0 21712 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_236
timestamp 1644511149
transform 1 0 22816 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_243
timestamp 1644511149
transform 1 0 23460 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_268
timestamp 1644511149
transform 1 0 25760 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_275
timestamp 1644511149
transform 1 0 26404 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_287
timestamp 1644511149
transform 1 0 27508 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_299
timestamp 1644511149
transform 1 0 28612 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1644511149
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_120
timestamp 1644511149
transform 1 0 12144 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_132
timestamp 1644511149
transform 1 0 13248 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_144
timestamp 1644511149
transform 1 0 14352 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_164
timestamp 1644511149
transform 1 0 16192 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_177
timestamp 1644511149
transform 1 0 17388 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_194
timestamp 1644511149
transform 1 0 18952 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_202
timestamp 1644511149
transform 1 0 19688 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_219
timestamp 1644511149
transform 1 0 21252 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_67_247
timestamp 1644511149
transform 1 0 23828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_269
timestamp 1644511149
transform 1 0 25852 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_276
timestamp 1644511149
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_115
timestamp 1644511149
transform 1 0 11684 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_123
timestamp 1644511149
transform 1 0 12420 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_127
timestamp 1644511149
transform 1 0 12788 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_134
timestamp 1644511149
transform 1 0 13432 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_149
timestamp 1644511149
transform 1 0 14812 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_158
timestamp 1644511149
transform 1 0 15640 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_178
timestamp 1644511149
transform 1 0 17480 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_187
timestamp 1644511149
transform 1 0 18308 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_200
timestamp 1644511149
transform 1 0 19504 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_212
timestamp 1644511149
transform 1 0 20608 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_221
timestamp 1644511149
transform 1 0 21436 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_225
timestamp 1644511149
transform 1 0 21804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_242
timestamp 1644511149
transform 1 0 23368 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_250
timestamp 1644511149
transform 1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_263
timestamp 1644511149
transform 1 0 25300 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_267
timestamp 1644511149
transform 1 0 25668 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_274
timestamp 1644511149
transform 1 0 26312 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_286
timestamp 1644511149
transform 1 0 27416 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_298
timestamp 1644511149
transform 1 0 28520 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_306
timestamp 1644511149
transform 1 0 29256 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_123
timestamp 1644511149
transform 1 0 12420 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_143
timestamp 1644511149
transform 1 0 14260 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_150
timestamp 1644511149
transform 1 0 14904 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_69_190
timestamp 1644511149
transform 1 0 18584 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_198
timestamp 1644511149
transform 1 0 19320 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_202
timestamp 1644511149
transform 1 0 19688 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_209
timestamp 1644511149
transform 1 0 20332 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_220
timestamp 1644511149
transform 1 0 21344 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_244
timestamp 1644511149
transform 1 0 23552 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_253
timestamp 1644511149
transform 1 0 24380 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1644511149
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1644511149
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_115
timestamp 1644511149
transform 1 0 11684 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_122
timestamp 1644511149
transform 1 0 12328 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_163
timestamp 1644511149
transform 1 0 16100 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_172
timestamp 1644511149
transform 1 0 16928 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_179
timestamp 1644511149
transform 1 0 17572 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_186
timestamp 1644511149
transform 1 0 18216 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_194
timestamp 1644511149
transform 1 0 18952 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_202
timestamp 1644511149
transform 1 0 19688 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_210
timestamp 1644511149
transform 1 0 20424 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_220
timestamp 1644511149
transform 1 0 21344 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_224
timestamp 1644511149
transform 1 0 21712 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1644511149
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1644511149
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1644511149
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1644511149
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1644511149
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1644511149
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1644511149
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_121
timestamp 1644511149
transform 1 0 12236 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_124
timestamp 1644511149
transform 1 0 12512 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_131
timestamp 1644511149
transform 1 0 13156 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_71_145
timestamp 1644511149
transform 1 0 14444 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_153
timestamp 1644511149
transform 1 0 15180 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_157
timestamp 1644511149
transform 1 0 15548 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_164
timestamp 1644511149
transform 1 0 16192 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_176
timestamp 1644511149
transform 1 0 17296 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_196
timestamp 1644511149
transform 1 0 19136 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_210
timestamp 1644511149
transform 1 0 20424 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_222
timestamp 1644511149
transform 1 0 21528 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_242
timestamp 1644511149
transform 1 0 23368 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_254
timestamp 1644511149
transform 1 0 24472 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_266
timestamp 1644511149
transform 1 0 25576 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_278
timestamp 1644511149
transform 1 0 26680 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1644511149
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1644511149
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_136
timestamp 1644511149
transform 1 0 13616 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_151
timestamp 1644511149
transform 1 0 14996 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_159
timestamp 1644511149
transform 1 0 15732 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_180
timestamp 1644511149
transform 1 0 17664 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_192
timestamp 1644511149
transform 1 0 18768 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_211
timestamp 1644511149
transform 1 0 20516 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_239
timestamp 1644511149
transform 1 0 23092 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_15
timestamp 1644511149
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_27
timestamp 1644511149
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_39
timestamp 1644511149
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1644511149
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_141
timestamp 1644511149
transform 1 0 14076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_150
timestamp 1644511149
transform 1 0 14904 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_162
timestamp 1644511149
transform 1 0 16008 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_179
timestamp 1644511149
transform 1 0 17572 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_186
timestamp 1644511149
transform 1 0 18216 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_194
timestamp 1644511149
transform 1 0 18952 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_203
timestamp 1644511149
transform 1 0 19780 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_215
timestamp 1644511149
transform 1 0 20884 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_243
timestamp 1644511149
transform 1 0 23460 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_252
timestamp 1644511149
transform 1 0 24288 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_264
timestamp 1644511149
transform 1 0 25392 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_276
timestamp 1644511149
transform 1 0 26496 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_129
timestamp 1644511149
transform 1 0 12972 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_136
timestamp 1644511149
transform 1 0 13616 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_149
timestamp 1644511149
transform 1 0 14812 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_203
timestamp 1644511149
transform 1 0 19780 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_219
timestamp 1644511149
transform 1 0 21252 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_228
timestamp 1644511149
transform 1 0 22080 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_237
timestamp 1644511149
transform 1 0 22908 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_249
timestamp 1644511149
transform 1 0 24012 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_258
timestamp 1644511149
transform 1 0 24840 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_262
timestamp 1644511149
transform 1 0 25208 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_274
timestamp 1644511149
transform 1 0 26312 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_286
timestamp 1644511149
transform 1 0 27416 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_298
timestamp 1644511149
transform 1 0 28520 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_306
timestamp 1644511149
transform 1 0 29256 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_15
timestamp 1644511149
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_27
timestamp 1644511149
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_39
timestamp 1644511149
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1644511149
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1644511149
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_142
timestamp 1644511149
transform 1 0 14168 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_154
timestamp 1644511149
transform 1 0 15272 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_158
timestamp 1644511149
transform 1 0 15640 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_164
timestamp 1644511149
transform 1 0 16192 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_185
timestamp 1644511149
transform 1 0 18124 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_197
timestamp 1644511149
transform 1 0 19228 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_203
timestamp 1644511149
transform 1 0 19780 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_209
timestamp 1644511149
transform 1 0 20332 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_221
timestamp 1644511149
transform 1 0 21436 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_245
timestamp 1644511149
transform 1 0 23644 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_251
timestamp 1644511149
transform 1 0 24196 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_258
timestamp 1644511149
transform 1 0 24840 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_270
timestamp 1644511149
transform 1 0 25944 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_278
timestamp 1644511149
transform 1 0 26680 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_146
timestamp 1644511149
transform 1 0 14536 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_174
timestamp 1644511149
transform 1 0 17112 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_188
timestamp 1644511149
transform 1 0 18400 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_213
timestamp 1644511149
transform 1 0 20700 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_231
timestamp 1644511149
transform 1 0 22356 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_235
timestamp 1644511149
transform 1 0 22724 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_242
timestamp 1644511149
transform 1 0 23368 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_250
timestamp 1644511149
transform 1 0 24104 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_289
timestamp 1644511149
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1644511149
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1644511149
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_144
timestamp 1644511149
transform 1 0 14352 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_164
timestamp 1644511149
transform 1 0 16192 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_188
timestamp 1644511149
transform 1 0 18400 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_200
timestamp 1644511149
transform 1 0 19504 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_219
timestamp 1644511149
transform 1 0 21252 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_77_243
timestamp 1644511149
transform 1 0 23460 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_250
timestamp 1644511149
transform 1 0 24104 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_262
timestamp 1644511149
transform 1 0 25208 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_274
timestamp 1644511149
transform 1 0 26312 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1644511149
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_181
timestamp 1644511149
transform 1 0 17756 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_192
timestamp 1644511149
transform 1 0 18768 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_208
timestamp 1644511149
transform 1 0 20240 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_216
timestamp 1644511149
transform 1 0 20976 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_222
timestamp 1644511149
transform 1 0 21528 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_234
timestamp 1644511149
transform 1 0 22632 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_248
timestamp 1644511149
transform 1 0 23920 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_289
timestamp 1644511149
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1644511149
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1644511149
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_15
timestamp 1644511149
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_27
timestamp 1644511149
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_39
timestamp 1644511149
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1644511149
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1644511149
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_131
timestamp 1644511149
transform 1 0 13156 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_145
timestamp 1644511149
transform 1 0 14444 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_157
timestamp 1644511149
transform 1 0 15548 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_165
timestamp 1644511149
transform 1 0 16284 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_175
timestamp 1644511149
transform 1 0 17204 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_199
timestamp 1644511149
transform 1 0 19412 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_208
timestamp 1644511149
transform 1 0 20240 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_214
timestamp 1644511149
transform 1 0 20792 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_220
timestamp 1644511149
transform 1 0 21344 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_229
timestamp 1644511149
transform 1 0 22172 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_235
timestamp 1644511149
transform 1 0 22724 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_243
timestamp 1644511149
transform 1 0 23460 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_255
timestamp 1644511149
transform 1 0 24564 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_267
timestamp 1644511149
transform 1 0 25668 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1644511149
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_309
timestamp 1644511149
transform 1 0 29532 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_314
timestamp 1644511149
transform 1 0 29992 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_326
timestamp 1644511149
transform 1 0 31096 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_334
timestamp 1644511149
transform 1 0 31832 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_337
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_349
timestamp 1644511149
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_361
timestamp 1644511149
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_373
timestamp 1644511149
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1644511149
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1644511149
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_15
timestamp 1644511149
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1644511149
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_41
timestamp 1644511149
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_53
timestamp 1644511149
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_65
timestamp 1644511149
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1644511149
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_109
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_80_122
timestamp 1644511149
transform 1 0 12328 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_135
timestamp 1644511149
transform 1 0 13524 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1644511149
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_141
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_150
timestamp 1644511149
transform 1 0 14904 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_159
timestamp 1644511149
transform 1 0 15732 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_168
timestamp 1644511149
transform 1 0 16560 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_177
timestamp 1644511149
transform 1 0 17388 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_184
timestamp 1644511149
transform 1 0 18032 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_209
timestamp 1644511149
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_221
timestamp 1644511149
transform 1 0 21436 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_232
timestamp 1644511149
transform 1 0 22448 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_244
timestamp 1644511149
transform 1 0 23552 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_265
timestamp 1644511149
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_277
timestamp 1644511149
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_289
timestamp 1644511149
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1644511149
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_333
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_345
timestamp 1644511149
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1644511149
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1644511149
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_395
timestamp 1644511149
transform 1 0 37444 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_403
timestamp 1644511149
transform 1 0 38180 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_15
timestamp 1644511149
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_27
timestamp 1644511149
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_39
timestamp 1644511149
transform 1 0 4692 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1644511149
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1644511149
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1644511149
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_119
timestamp 1644511149
transform 1 0 12052 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_123
timestamp 1644511149
transform 1 0 12420 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_130
timestamp 1644511149
transform 1 0 13064 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_139
timestamp 1644511149
transform 1 0 13892 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_146
timestamp 1644511149
transform 1 0 14536 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_81_157
timestamp 1644511149
transform 1 0 15548 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_164
timestamp 1644511149
transform 1 0 16192 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_174
timestamp 1644511149
transform 1 0 17112 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_178
timestamp 1644511149
transform 1 0 17480 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_183
timestamp 1644511149
transform 1 0 17940 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_81_192
timestamp 1644511149
transform 1 0 18768 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_203
timestamp 1644511149
transform 1 0 19780 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_215
timestamp 1644511149
transform 1 0 20884 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_219
timestamp 1644511149
transform 1 0 21252 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1644511149
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_229
timestamp 1644511149
transform 1 0 22172 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_241
timestamp 1644511149
transform 1 0 23276 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_81_250
timestamp 1644511149
transform 1 0 24104 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_262
timestamp 1644511149
transform 1 0 25208 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_274
timestamp 1644511149
transform 1 0 26312 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_81_285
timestamp 1644511149
transform 1 0 27324 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_297
timestamp 1644511149
transform 1 0 28428 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_309
timestamp 1644511149
transform 1 0 29532 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_320
timestamp 1644511149
transform 1 0 30544 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_332
timestamp 1644511149
transform 1 0 31648 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_340
timestamp 1644511149
transform 1 0 32384 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_81_349
timestamp 1644511149
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_361
timestamp 1644511149
transform 1 0 34316 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_368
timestamp 1644511149
transform 1 0 34960 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_380
timestamp 1644511149
transform 1 0 36064 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_403
timestamp 1644511149
transform 1 0 38180 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_7
timestamp 1644511149
transform 1 0 1748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_15
timestamp 1644511149
transform 1 0 2484 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_23
timestamp 1644511149
transform 1 0 3220 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_33
timestamp 1644511149
transform 1 0 4140 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_41
timestamp 1644511149
transform 1 0 4876 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_49
timestamp 1644511149
transform 1 0 5612 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_55
timestamp 1644511149
transform 1 0 6164 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_61
timestamp 1644511149
transform 1 0 6716 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_69
timestamp 1644511149
transform 1 0 7452 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_73
timestamp 1644511149
transform 1 0 7820 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_78
timestamp 1644511149
transform 1 0 8280 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_89
timestamp 1644511149
transform 1 0 9292 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_97
timestamp 1644511149
transform 1 0 10028 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_105
timestamp 1644511149
transform 1 0 10764 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_111
timestamp 1644511149
transform 1 0 11316 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_117
timestamp 1644511149
transform 1 0 11868 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_125
timestamp 1644511149
transform 1 0 12604 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1644511149
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1644511149
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_145
timestamp 1644511149
transform 1 0 14444 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_153
timestamp 1644511149
transform 1 0 15180 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_161
timestamp 1644511149
transform 1 0 15916 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_167
timestamp 1644511149
transform 1 0 16468 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_173
timestamp 1644511149
transform 1 0 17020 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_181
timestamp 1644511149
transform 1 0 17756 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1644511149
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1644511149
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_201
timestamp 1644511149
transform 1 0 19596 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_209
timestamp 1644511149
transform 1 0 20332 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_217
timestamp 1644511149
transform 1 0 21068 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_223
timestamp 1644511149
transform 1 0 21620 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_82_225
timestamp 1644511149
transform 1 0 21804 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_232
timestamp 1644511149
transform 1 0 22448 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_236
timestamp 1644511149
transform 1 0 22816 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_241
timestamp 1644511149
transform 1 0 23276 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_249
timestamp 1644511149
transform 1 0 24012 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_257
timestamp 1644511149
transform 1 0 24748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_265
timestamp 1644511149
transform 1 0 25484 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_273
timestamp 1644511149
transform 1 0 26220 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_279
timestamp 1644511149
transform 1 0 26772 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_281
timestamp 1644511149
transform 1 0 26956 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_289
timestamp 1644511149
transform 1 0 27692 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_297
timestamp 1644511149
transform 1 0 28428 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_305
timestamp 1644511149
transform 1 0 29164 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_319
timestamp 1644511149
transform 1 0 30452 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_327
timestamp 1644511149
transform 1 0 31188 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_331
timestamp 1644511149
transform 1 0 31556 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_335
timestamp 1644511149
transform 1 0 31924 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_347
timestamp 1644511149
transform 1 0 33028 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_359
timestamp 1644511149
transform 1 0 34132 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1644511149
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_369
timestamp 1644511149
transform 1 0 35052 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_374
timestamp 1644511149
transform 1 0 35512 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_388
timestamp 1644511149
transform 1 0 36800 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_403
timestamp 1644511149
transform 1 0 38180 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 38824 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 38824 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 38824 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 38824 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 38824 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 38824 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 38824 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 38824 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 38824 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 38824 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 38824 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 38824 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 38824 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 38824 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 38824 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 38824 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 38824 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 38824 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _0968_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14996 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0969_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0970_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26128 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0971_
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0972_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0973_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23000 0 1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0974_
timestamp 1644511149
transform 1 0 28336 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0975_
timestamp 1644511149
transform 1 0 28428 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0976_
timestamp 1644511149
transform 1 0 28244 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0977_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27508 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0978_
timestamp 1644511149
transform 1 0 27784 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0979_
timestamp 1644511149
transform 1 0 28428 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0980_
timestamp 1644511149
transform 1 0 27508 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0981_
timestamp 1644511149
transform 1 0 27324 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0982_
timestamp 1644511149
transform 1 0 24472 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0983_
timestamp 1644511149
transform 1 0 25944 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0984_
timestamp 1644511149
transform 1 0 25024 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0985_
timestamp 1644511149
transform 1 0 24656 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0986_
timestamp 1644511149
transform 1 0 23184 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0987_
timestamp 1644511149
transform 1 0 23000 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0988_
timestamp 1644511149
transform 1 0 23000 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0989_
timestamp 1644511149
transform 1 0 22540 0 -1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0990_
timestamp 1644511149
transform 1 0 18308 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0991_
timestamp 1644511149
transform 1 0 19320 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0992_
timestamp 1644511149
transform 1 0 18768 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0993_
timestamp 1644511149
transform 1 0 19320 0 1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0994_
timestamp 1644511149
transform 1 0 18676 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0995_
timestamp 1644511149
transform 1 0 17296 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0996_
timestamp 1644511149
transform 1 0 17020 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0997_
timestamp 1644511149
transform 1 0 17480 0 1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0998_
timestamp 1644511149
transform 1 0 13156 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0999_
timestamp 1644511149
transform 1 0 12512 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1000_
timestamp 1644511149
transform 1 0 11776 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1001_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1002_
timestamp 1644511149
transform 1 0 25116 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1003_
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1004_
timestamp 1644511149
transform 1 0 24748 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1005_
timestamp 1644511149
transform 1 0 24748 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1006_
timestamp 1644511149
transform 1 0 31188 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1007_
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1008_
timestamp 1644511149
transform 1 0 29900 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1009_
timestamp 1644511149
transform 1 0 29624 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1010_
timestamp 1644511149
transform 1 0 30912 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1011_
timestamp 1644511149
transform 1 0 31096 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1012_
timestamp 1644511149
transform 1 0 29256 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1013_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1014_
timestamp 1644511149
transform 1 0 23644 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1015_
timestamp 1644511149
transform 1 0 24104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1016_
timestamp 1644511149
transform 1 0 23368 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1017_
timestamp 1644511149
transform 1 0 23092 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1018_
timestamp 1644511149
transform 1 0 20700 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1019_
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1020_
timestamp 1644511149
transform 1 0 21344 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1021_
timestamp 1644511149
transform 1 0 21160 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1022_
timestamp 1644511149
transform 1 0 17940 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1023_
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1024_
timestamp 1644511149
transform 1 0 18216 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1025_
timestamp 1644511149
transform 1 0 17848 0 1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1026_
timestamp 1644511149
transform 1 0 15824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1027_
timestamp 1644511149
transform 1 0 13340 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1028_
timestamp 1644511149
transform 1 0 12972 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1029_
timestamp 1644511149
transform 1 0 13524 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1030_
timestamp 1644511149
transform 1 0 11776 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1031_
timestamp 1644511149
transform 1 0 12328 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1032_
timestamp 1644511149
transform 1 0 11592 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1033_
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1034_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22264 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1035_
timestamp 1644511149
transform 1 0 23828 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1036_
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1037_
timestamp 1644511149
transform 1 0 24564 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1038_
timestamp 1644511149
transform 1 0 23828 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1644511149
transform 1 0 23920 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1040_
timestamp 1644511149
transform 1 0 22908 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1644511149
transform 1 0 23828 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1042_
timestamp 1644511149
transform 1 0 20884 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1043_
timestamp 1644511149
transform 1 0 22172 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1044_
timestamp 1644511149
transform 1 0 19780 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1045_
timestamp 1644511149
transform 1 0 20976 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1046_
timestamp 1644511149
transform 1 0 17940 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1047_
timestamp 1644511149
transform 1 0 19136 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1048_
timestamp 1644511149
transform 1 0 14444 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1049_
timestamp 1644511149
transform 1 0 19504 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1050_
timestamp 1644511149
transform 1 0 17296 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1051_
timestamp 1644511149
transform 1 0 18492 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1052_
timestamp 1644511149
transform 1 0 15272 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1053_
timestamp 1644511149
transform 1 0 17664 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1054_
timestamp 1644511149
transform 1 0 16928 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1055_
timestamp 1644511149
transform 1 0 17756 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1056_
timestamp 1644511149
transform 1 0 16100 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1057_
timestamp 1644511149
transform 1 0 15916 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1058_
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1059_
timestamp 1644511149
transform 1 0 15272 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1060_
timestamp 1644511149
transform 1 0 13064 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1061_
timestamp 1644511149
transform 1 0 14260 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1062_
timestamp 1644511149
transform 1 0 13432 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1063_
timestamp 1644511149
transform 1 0 12788 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1064_
timestamp 1644511149
transform 1 0 11868 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1065_
timestamp 1644511149
transform 1 0 12144 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1066_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17940 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1067_
timestamp 1644511149
transform 1 0 19596 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1068_
timestamp 1644511149
transform 1 0 19596 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1069_
timestamp 1644511149
transform 1 0 15456 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _1070_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1071_
timestamp 1644511149
transform 1 0 16100 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1072_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32384 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1073_
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1074_
timestamp 1644511149
transform 1 0 28520 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1075_
timestamp 1644511149
transform 1 0 24472 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1076_
timestamp 1644511149
transform 1 0 29348 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1077_
timestamp 1644511149
transform 1 0 18032 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1078_
timestamp 1644511149
transform 1 0 18124 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1079_
timestamp 1644511149
transform 1 0 15364 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1080_
timestamp 1644511149
transform 1 0 18952 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1081_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16192 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1082_
timestamp 1644511149
transform 1 0 15456 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1083_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14628 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1084_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_4  _1085_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14628 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1086_
timestamp 1644511149
transform 1 0 15180 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1087_
timestamp 1644511149
transform 1 0 14352 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1088_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14904 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_4  _1089_
timestamp 1644511149
transform 1 0 14720 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1090_
timestamp 1644511149
transform 1 0 14904 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__or3_4  _1091_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _1092_
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1093_
timestamp 1644511149
transform 1 0 16192 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or2_2  _1094_
timestamp 1644511149
transform 1 0 15272 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1095_
timestamp 1644511149
transform 1 0 13984 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _1096_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16836 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1097_
timestamp 1644511149
transform 1 0 15824 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _1098_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17204 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  _1099_
timestamp 1644511149
transform 1 0 22632 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1100_
timestamp 1644511149
transform 1 0 28796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1101_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11960 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1102_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12144 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_2  _1103_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16928 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1104_
timestamp 1644511149
transform 1 0 17388 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1105_
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1106_
timestamp 1644511149
transform 1 0 11684 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1107_
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1108_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19964 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1109_
timestamp 1644511149
transform 1 0 16008 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1110_
timestamp 1644511149
transform 1 0 16836 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _1111_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17848 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _1112_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1113_
timestamp 1644511149
transform 1 0 17296 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1114_
timestamp 1644511149
transform 1 0 16376 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1115_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11408 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1116_
timestamp 1644511149
transform 1 0 17664 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1117_
timestamp 1644511149
transform 1 0 18400 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1118_
timestamp 1644511149
transform 1 0 23276 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1119_
timestamp 1644511149
transform 1 0 16376 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1120_
timestamp 1644511149
transform 1 0 16744 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1121_
timestamp 1644511149
transform 1 0 16008 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1122_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15548 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _1123_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15180 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1124_
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1125_
timestamp 1644511149
transform 1 0 25024 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1126_
timestamp 1644511149
transform 1 0 23000 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1127_
timestamp 1644511149
transform 1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1128_
timestamp 1644511149
transform 1 0 14628 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1129_
timestamp 1644511149
transform 1 0 12052 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1130_
timestamp 1644511149
transform 1 0 12052 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1131_
timestamp 1644511149
transform 1 0 11592 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1132_
timestamp 1644511149
transform 1 0 10764 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1133_
timestamp 1644511149
transform 1 0 17940 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1134_
timestamp 1644511149
transform 1 0 17572 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1135_
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1136_
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1137_
timestamp 1644511149
transform 1 0 19228 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__a32o_1  _1138_
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1139_
timestamp 1644511149
transform 1 0 16192 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1140_
timestamp 1644511149
transform 1 0 21712 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1141_
timestamp 1644511149
transform 1 0 21712 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1142_
timestamp 1644511149
transform 1 0 16652 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1143_
timestamp 1644511149
transform 1 0 15456 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1144_
timestamp 1644511149
transform 1 0 20148 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1145_
timestamp 1644511149
transform 1 0 14720 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1146_
timestamp 1644511149
transform 1 0 14628 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1147_
timestamp 1644511149
transform 1 0 10580 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1148_
timestamp 1644511149
transform 1 0 10672 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1149_
timestamp 1644511149
transform 1 0 15640 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1150_
timestamp 1644511149
transform 1 0 17848 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1151_
timestamp 1644511149
transform 1 0 16744 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1152_
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1153_
timestamp 1644511149
transform 1 0 17112 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1154_
timestamp 1644511149
transform 1 0 16560 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1155_
timestamp 1644511149
transform 1 0 13616 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1156_
timestamp 1644511149
transform 1 0 13616 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1157_
timestamp 1644511149
transform 1 0 12972 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1158_
timestamp 1644511149
transform 1 0 12880 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1159_
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1160_
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _1161_
timestamp 1644511149
transform 1 0 15916 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1162_
timestamp 1644511149
transform 1 0 13340 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1163_
timestamp 1644511149
transform 1 0 15916 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1164_
timestamp 1644511149
transform 1 0 14352 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1165_
timestamp 1644511149
transform 1 0 15272 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1166_
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1167_
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1168_
timestamp 1644511149
transform 1 0 12880 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1169_
timestamp 1644511149
transform 1 0 17848 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1170_
timestamp 1644511149
transform 1 0 18216 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _1171_
timestamp 1644511149
transform 1 0 17572 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1172_
timestamp 1644511149
transform 1 0 18584 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1173_
timestamp 1644511149
transform 1 0 17112 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1174_
timestamp 1644511149
transform 1 0 16560 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1175_
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1176_
timestamp 1644511149
transform 1 0 19780 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__a32o_1  _1177_
timestamp 1644511149
transform 1 0 18676 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1178_
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1179_
timestamp 1644511149
transform 1 0 23000 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1180_
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1181_
timestamp 1644511149
transform 1 0 18124 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1182_
timestamp 1644511149
transform 1 0 18032 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1183_
timestamp 1644511149
transform 1 0 19872 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1184_
timestamp 1644511149
transform 1 0 20424 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1185_
timestamp 1644511149
transform 1 0 18676 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1186_
timestamp 1644511149
transform 1 0 17940 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1187_
timestamp 1644511149
transform 1 0 19688 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1188_
timestamp 1644511149
transform 1 0 20884 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _1189_
timestamp 1644511149
transform 1 0 20056 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1190_
timestamp 1644511149
transform 1 0 19596 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1191_
timestamp 1644511149
transform 1 0 19412 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1192_
timestamp 1644511149
transform 1 0 20516 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1193_
timestamp 1644511149
transform 1 0 21620 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1194_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1195_
timestamp 1644511149
transform 1 0 20056 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1196_
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1197_
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _1198_
timestamp 1644511149
transform 1 0 20700 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1199_
timestamp 1644511149
transform 1 0 22172 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1200_
timestamp 1644511149
transform 1 0 21068 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1201_
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1202_
timestamp 1644511149
transform 1 0 20792 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1203_
timestamp 1644511149
transform 1 0 18032 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1204_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19688 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1205_
timestamp 1644511149
transform 1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1206_
timestamp 1644511149
transform 1 0 20608 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1207_
timestamp 1644511149
transform 1 0 19688 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1208_
timestamp 1644511149
transform 1 0 20608 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1209_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18952 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1210_
timestamp 1644511149
transform 1 0 27508 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1211_
timestamp 1644511149
transform 1 0 20976 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1212_
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1213_
timestamp 1644511149
transform 1 0 23552 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _1214_
timestamp 1644511149
transform 1 0 17112 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  _1215_
timestamp 1644511149
transform 1 0 26220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1216_
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1217_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1218_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1219_
timestamp 1644511149
transform 1 0 23644 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1220_
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1221_
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1222_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1223_
timestamp 1644511149
transform 1 0 23644 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1224_
timestamp 1644511149
transform 1 0 24472 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1225_
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1226_
timestamp 1644511149
transform 1 0 26220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1227_
timestamp 1644511149
transform 1 0 24932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1228_
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1229_
timestamp 1644511149
transform 1 0 26036 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1230_
timestamp 1644511149
transform 1 0 25760 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1231_
timestamp 1644511149
transform 1 0 25668 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1232_
timestamp 1644511149
transform 1 0 25392 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1233_
timestamp 1644511149
transform 1 0 27140 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1234_
timestamp 1644511149
transform 1 0 26312 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1235_
timestamp 1644511149
transform 1 0 26956 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1236_
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1237_
timestamp 1644511149
transform 1 0 29808 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1238_
timestamp 1644511149
transform 1 0 30452 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1239_
timestamp 1644511149
transform 1 0 29808 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1240_
timestamp 1644511149
transform 1 0 29716 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1241_
timestamp 1644511149
transform 1 0 25760 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1242_
timestamp 1644511149
transform 1 0 26956 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1243_
timestamp 1644511149
transform 1 0 27784 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1244_
timestamp 1644511149
transform 1 0 27968 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1245_
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1246_
timestamp 1644511149
transform 1 0 30084 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1247_
timestamp 1644511149
transform 1 0 30360 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1248_
timestamp 1644511149
transform 1 0 30636 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1249_
timestamp 1644511149
transform 1 0 31372 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1250_
timestamp 1644511149
transform 1 0 27876 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1251_
timestamp 1644511149
transform 1 0 27968 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1252_
timestamp 1644511149
transform 1 0 28244 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1253_
timestamp 1644511149
transform 1 0 30360 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1254_
timestamp 1644511149
transform 1 0 32476 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1255_
timestamp 1644511149
transform 1 0 32568 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1256_
timestamp 1644511149
transform 1 0 33028 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1257_
timestamp 1644511149
transform 1 0 28520 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1258_
timestamp 1644511149
transform 1 0 28704 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1259_
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1260_
timestamp 1644511149
transform 1 0 30360 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1261_
timestamp 1644511149
transform 1 0 33764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1262_
timestamp 1644511149
transform 1 0 32936 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1263_
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1264_
timestamp 1644511149
transform 1 0 27784 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1265_
timestamp 1644511149
transform 1 0 28336 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1266_
timestamp 1644511149
transform 1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1267_
timestamp 1644511149
transform 1 0 25668 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1268_
timestamp 1644511149
transform 1 0 33672 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1269_
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1270_
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1271_
timestamp 1644511149
transform 1 0 25760 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _1272_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1273_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28336 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1274_
timestamp 1644511149
transform 1 0 24564 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1275_
timestamp 1644511149
transform 1 0 32292 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1276_
timestamp 1644511149
transform 1 0 33028 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1277_
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1278_
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1279_
timestamp 1644511149
transform 1 0 12420 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1280_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13064 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1281_
timestamp 1644511149
transform 1 0 11684 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1282_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11684 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1283_
timestamp 1644511149
transform 1 0 11408 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1284_
timestamp 1644511149
transform 1 0 14720 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1285_
timestamp 1644511149
transform 1 0 13984 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1286_
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1287_
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1288_
timestamp 1644511149
transform 1 0 19136 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1289_
timestamp 1644511149
transform 1 0 20516 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1290_
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1291_
timestamp 1644511149
transform 1 0 11592 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1292_
timestamp 1644511149
transform 1 0 22080 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1293_
timestamp 1644511149
transform 1 0 22632 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1294_
timestamp 1644511149
transform 1 0 21896 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1295_
timestamp 1644511149
transform 1 0 22264 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1296_
timestamp 1644511149
transform 1 0 23460 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1297_
timestamp 1644511149
transform 1 0 24380 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1298_
timestamp 1644511149
transform 1 0 23276 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1299_
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1300_
timestamp 1644511149
transform 1 0 13340 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1301_
timestamp 1644511149
transform 1 0 30820 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1302_
timestamp 1644511149
transform 1 0 30728 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1303_
timestamp 1644511149
transform 1 0 30084 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1304_
timestamp 1644511149
transform 1 0 30544 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1305_
timestamp 1644511149
transform 1 0 30360 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1306_
timestamp 1644511149
transform 1 0 30176 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1307_
timestamp 1644511149
transform 1 0 30176 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1308_
timestamp 1644511149
transform 1 0 31188 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1309_
timestamp 1644511149
transform 1 0 25852 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1310_
timestamp 1644511149
transform 1 0 26128 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1311_
timestamp 1644511149
transform 1 0 25116 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1312_
timestamp 1644511149
transform 1 0 26220 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1313_
timestamp 1644511149
transform 1 0 12696 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1314_
timestamp 1644511149
transform 1 0 13156 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1315_
timestamp 1644511149
transform 1 0 12696 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1316_
timestamp 1644511149
transform 1 0 14628 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1317_
timestamp 1644511149
transform 1 0 15732 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1318_
timestamp 1644511149
transform 1 0 17940 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1319_
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1320_
timestamp 1644511149
transform 1 0 17940 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1321_
timestamp 1644511149
transform 1 0 18952 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1322_
timestamp 1644511149
transform 1 0 19872 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1323_
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1324_
timestamp 1644511149
transform 1 0 19412 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1325_
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1326_
timestamp 1644511149
transform 1 0 23920 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1327_
timestamp 1644511149
transform 1 0 23644 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1328_
timestamp 1644511149
transform 1 0 23276 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1329_
timestamp 1644511149
transform 1 0 24288 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1330_
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1331_
timestamp 1644511149
transform 1 0 25668 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1332_
timestamp 1644511149
transform 1 0 25484 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1333_
timestamp 1644511149
transform 1 0 26312 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1334_
timestamp 1644511149
transform 1 0 27876 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1335_
timestamp 1644511149
transform 1 0 28796 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1336_
timestamp 1644511149
transform 1 0 27784 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1337_
timestamp 1644511149
transform 1 0 27876 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1338_
timestamp 1644511149
transform 1 0 29164 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1339_
timestamp 1644511149
transform 1 0 28704 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1340_
timestamp 1644511149
transform 1 0 28244 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1341_
timestamp 1644511149
transform 1 0 27600 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1342_
timestamp 1644511149
transform 1 0 18400 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1343_
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1344_
timestamp 1644511149
transform 1 0 24656 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1345_
timestamp 1644511149
transform 1 0 23828 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1346_
timestamp 1644511149
transform 1 0 17480 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1347_
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1348_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18124 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _1349_
timestamp 1644511149
transform 1 0 16928 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1350_
timestamp 1644511149
transform 1 0 20792 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1351_
timestamp 1644511149
transform 1 0 20056 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1352_
timestamp 1644511149
transform 1 0 9292 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1353_
timestamp 1644511149
transform 1 0 10396 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1354_
timestamp 1644511149
transform 1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1355_
timestamp 1644511149
transform 1 0 31556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1356_
timestamp 1644511149
transform 1 0 31924 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1357_
timestamp 1644511149
transform 1 0 32936 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1358_
timestamp 1644511149
transform 1 0 9292 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1359_
timestamp 1644511149
transform 1 0 7728 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1360_
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1361_
timestamp 1644511149
transform 1 0 5428 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1362_
timestamp 1644511149
transform 1 0 4784 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1363_
timestamp 1644511149
transform 1 0 31096 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1364_
timestamp 1644511149
transform 1 0 32936 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1365_
timestamp 1644511149
transform 1 0 7452 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1366_
timestamp 1644511149
transform 1 0 5336 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1367_
timestamp 1644511149
transform 1 0 4232 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1368_
timestamp 1644511149
transform 1 0 32108 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1369_
timestamp 1644511149
transform 1 0 33764 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1370_
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1371_
timestamp 1644511149
transform 1 0 2852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1372_
timestamp 1644511149
transform 1 0 32108 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1373_
timestamp 1644511149
transform 1 0 33764 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1374_
timestamp 1644511149
transform 1 0 4600 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1375_
timestamp 1644511149
transform 1 0 4876 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1376_
timestamp 1644511149
transform 1 0 32568 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1377_
timestamp 1644511149
transform 1 0 34500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1378_
timestamp 1644511149
transform 1 0 4508 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1379_
timestamp 1644511149
transform 1 0 4324 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1380_
timestamp 1644511149
transform 1 0 31556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1381_
timestamp 1644511149
transform 1 0 31188 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1382_
timestamp 1644511149
transform 1 0 33580 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1383_
timestamp 1644511149
transform 1 0 6716 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1384_
timestamp 1644511149
transform 1 0 6440 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1385_
timestamp 1644511149
transform 1 0 5612 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1386_
timestamp 1644511149
transform 1 0 30268 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1387_
timestamp 1644511149
transform 1 0 33580 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1388_
timestamp 1644511149
transform 1 0 8464 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1389_
timestamp 1644511149
transform 1 0 7360 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1390_
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1391_
timestamp 1644511149
transform 1 0 32936 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1392_
timestamp 1644511149
transform 1 0 32752 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1393_
timestamp 1644511149
transform 1 0 7360 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1394_
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1395_
timestamp 1644511149
transform 1 0 32936 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1396_
timestamp 1644511149
transform 1 0 33396 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1397_
timestamp 1644511149
transform 1 0 7360 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1398_
timestamp 1644511149
transform 1 0 10396 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1399_
timestamp 1644511149
transform 1 0 33396 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1400_
timestamp 1644511149
transform 1 0 32016 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1401_
timestamp 1644511149
transform 1 0 7636 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1402_
timestamp 1644511149
transform 1 0 8096 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1403_
timestamp 1644511149
transform 1 0 30912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1404_
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1405_
timestamp 1644511149
transform 1 0 29624 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1406_
timestamp 1644511149
transform 1 0 7360 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1407_
timestamp 1644511149
transform 1 0 6532 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1408_
timestamp 1644511149
transform 1 0 6256 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1409_
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1410_
timestamp 1644511149
transform 1 0 36340 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1411_
timestamp 1644511149
transform 1 0 8280 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1412_
timestamp 1644511149
transform 1 0 6900 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1413_
timestamp 1644511149
transform 1 0 6716 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1414_
timestamp 1644511149
transform 1 0 31280 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1415_
timestamp 1644511149
transform 1 0 36340 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1416_
timestamp 1644511149
transform 1 0 8004 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1417_
timestamp 1644511149
transform 1 0 6716 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1418_
timestamp 1644511149
transform 1 0 30360 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1419_
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1420_
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1421_
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1422_
timestamp 1644511149
transform 1 0 32568 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1423_
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1424_
timestamp 1644511149
transform 1 0 5152 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1425_
timestamp 1644511149
transform 1 0 4508 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1426_
timestamp 1644511149
transform 1 0 30544 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1427_
timestamp 1644511149
transform 1 0 30268 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1428_
timestamp 1644511149
transform 1 0 6624 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _1429_
timestamp 1644511149
transform 1 0 16928 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1430_
timestamp 1644511149
transform 1 0 10488 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1431_
timestamp 1644511149
transform 1 0 10488 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1432_
timestamp 1644511149
transform 1 0 7728 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1433_
timestamp 1644511149
transform 1 0 7728 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1434_
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1435_
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1436_
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1437_
timestamp 1644511149
transform 1 0 7176 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1438_
timestamp 1644511149
transform 1 0 7728 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1439_
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1440_
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1441_
timestamp 1644511149
transform 1 0 8004 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1442_
timestamp 1644511149
transform 1 0 9752 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1443_
timestamp 1644511149
transform 1 0 7728 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1444_
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1445_
timestamp 1644511149
transform 1 0 5612 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1446_
timestamp 1644511149
transform 1 0 7452 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1447_
timestamp 1644511149
transform 1 0 4784 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1448_
timestamp 1644511149
transform 1 0 5428 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1449_
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1450_
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1451_
timestamp 1644511149
transform 1 0 4784 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1452_
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1453_
timestamp 1644511149
transform 1 0 6256 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1454_
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1455_
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1456_
timestamp 1644511149
transform 1 0 7176 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1457_
timestamp 1644511149
transform 1 0 7728 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1458_
timestamp 1644511149
transform 1 0 7728 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1459_
timestamp 1644511149
transform 1 0 8648 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1460_
timestamp 1644511149
transform 1 0 6164 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1461_
timestamp 1644511149
transform 1 0 9292 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1462_
timestamp 1644511149
transform 1 0 7728 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1463_
timestamp 1644511149
transform 1 0 7820 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1464_
timestamp 1644511149
transform 1 0 5428 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1465_
timestamp 1644511149
transform 1 0 6256 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1466_
timestamp 1644511149
transform 1 0 9752 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1467_
timestamp 1644511149
transform 1 0 7728 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1468_
timestamp 1644511149
transform 1 0 8464 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1469_
timestamp 1644511149
transform 1 0 5428 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1470_
timestamp 1644511149
transform 1 0 6256 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1471_
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1472_
timestamp 1644511149
transform 1 0 5520 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1473_
timestamp 1644511149
transform 1 0 7176 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1474_
timestamp 1644511149
transform 1 0 5612 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1475_
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1476_
timestamp 1644511149
transform 1 0 5428 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1477_
timestamp 1644511149
transform 1 0 8188 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1478_
timestamp 1644511149
transform 1 0 9568 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1479_
timestamp 1644511149
transform 1 0 12604 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1480_
timestamp 1644511149
transform 1 0 11868 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1481_
timestamp 1644511149
transform 1 0 9844 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1482_
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1483_
timestamp 1644511149
transform 1 0 9936 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1484_
timestamp 1644511149
transform 1 0 7820 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1485_
timestamp 1644511149
transform 1 0 5612 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1486_
timestamp 1644511149
transform 1 0 10672 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1487_
timestamp 1644511149
transform 1 0 9568 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1488_
timestamp 1644511149
transform 1 0 6992 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1489_
timestamp 1644511149
transform 1 0 7176 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1490_
timestamp 1644511149
transform 1 0 11224 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1491_
timestamp 1644511149
transform 1 0 10396 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1492_
timestamp 1644511149
transform 1 0 10028 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1493_
timestamp 1644511149
transform 1 0 7176 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1494_
timestamp 1644511149
transform 1 0 6900 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1495_
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1496_
timestamp 1644511149
transform 1 0 11316 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1497_
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1498_
timestamp 1644511149
transform 1 0 7820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1499_
timestamp 1644511149
transform 1 0 12604 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1500_
timestamp 1644511149
transform 1 0 12328 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1501_
timestamp 1644511149
transform 1 0 9016 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1502_
timestamp 1644511149
transform 1 0 7912 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1503_
timestamp 1644511149
transform 1 0 12696 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1504_
timestamp 1644511149
transform 1 0 11776 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1505_
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1506_
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1507_
timestamp 1644511149
transform 1 0 8464 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1508_
timestamp 1644511149
transform 1 0 12512 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _1509_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2852 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1510_
timestamp 1644511149
transform 1 0 16100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1511_
timestamp 1644511149
transform 1 0 23000 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1512_
timestamp 1644511149
transform 1 0 23184 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1513_
timestamp 1644511149
transform 1 0 13340 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1514_
timestamp 1644511149
transform 1 0 23184 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _1515_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10764 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1516_
timestamp 1644511149
transform 1 0 12328 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1517_
timestamp 1644511149
transform 1 0 19688 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1518_
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1519_
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1520_
timestamp 1644511149
transform 1 0 19504 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1521_
timestamp 1644511149
transform 1 0 17572 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1522_
timestamp 1644511149
transform 1 0 18032 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1523_
timestamp 1644511149
transform 1 0 18124 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1524_
timestamp 1644511149
transform 1 0 15364 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1525_
timestamp 1644511149
transform 1 0 8188 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1526_
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1527_
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1528_
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1529_
timestamp 1644511149
transform 1 0 23736 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1530_
timestamp 1644511149
transform 1 0 25392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1531_
timestamp 1644511149
transform 1 0 15456 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_1  _1532_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10028 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1533_
timestamp 1644511149
transform 1 0 10212 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1534_
timestamp 1644511149
transform 1 0 8004 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1535_
timestamp 1644511149
transform 1 0 9016 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1536_
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1537_
timestamp 1644511149
transform 1 0 10580 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1538_
timestamp 1644511149
transform 1 0 9936 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1539_
timestamp 1644511149
transform 1 0 17020 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1540_
timestamp 1644511149
transform 1 0 9660 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1541_
timestamp 1644511149
transform 1 0 10672 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1542_
timestamp 1644511149
transform 1 0 10120 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1543_
timestamp 1644511149
transform 1 0 10120 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1544_
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1545_
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1546_
timestamp 1644511149
transform 1 0 11592 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1547_
timestamp 1644511149
transform 1 0 11776 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1548_
timestamp 1644511149
transform 1 0 12236 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1549_
timestamp 1644511149
transform 1 0 13064 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1550_
timestamp 1644511149
transform 1 0 19596 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1551_
timestamp 1644511149
transform 1 0 20976 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1552_
timestamp 1644511149
transform 1 0 14444 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1553_
timestamp 1644511149
transform 1 0 14628 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1554_
timestamp 1644511149
transform 1 0 15456 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1555_
timestamp 1644511149
transform 1 0 14904 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_1  _1556_
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1557_
timestamp 1644511149
transform 1 0 12788 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1558_
timestamp 1644511149
transform 1 0 19596 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1559_
timestamp 1644511149
transform 1 0 17480 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1560_
timestamp 1644511149
transform 1 0 18308 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1561_
timestamp 1644511149
transform 1 0 17480 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1562_
timestamp 1644511149
transform 1 0 23000 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1563_
timestamp 1644511149
transform 1 0 23920 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_1  _1564_
timestamp 1644511149
transform 1 0 19136 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1565_
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1566_
timestamp 1644511149
transform 1 0 18492 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1567_
timestamp 1644511149
transform 1 0 18308 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1568_
timestamp 1644511149
transform 1 0 18952 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1569_
timestamp 1644511149
transform 1 0 19596 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1570_
timestamp 1644511149
transform 1 0 20608 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1571_
timestamp 1644511149
transform 1 0 20148 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1572_
timestamp 1644511149
transform 1 0 20608 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1573_
timestamp 1644511149
transform 1 0 21160 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1574_
timestamp 1644511149
transform 1 0 20884 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1575_
timestamp 1644511149
transform 1 0 21160 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1576_
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1577_
timestamp 1644511149
transform 1 0 21988 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1578_
timestamp 1644511149
transform 1 0 22264 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1579_
timestamp 1644511149
transform 1 0 21620 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1580_
timestamp 1644511149
transform 1 0 22724 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1581_
timestamp 1644511149
transform 1 0 23552 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1582_
timestamp 1644511149
transform 1 0 23000 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1583_
timestamp 1644511149
transform 1 0 24380 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1584_
timestamp 1644511149
transform 1 0 24288 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1585_
timestamp 1644511149
transform 1 0 25116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1586_
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_1  _1587_
timestamp 1644511149
transform 1 0 24748 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1588_
timestamp 1644511149
transform 1 0 25576 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1589_
timestamp 1644511149
transform 1 0 25024 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1590_
timestamp 1644511149
transform 1 0 26496 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1591_
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1592_
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1593_
timestamp 1644511149
transform 1 0 24748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1594_
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__o22ai_1  _1595_
timestamp 1644511149
transform 1 0 27508 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1596_
timestamp 1644511149
transform 1 0 27416 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1597_
timestamp 1644511149
transform 1 0 28428 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1598_
timestamp 1644511149
transform 1 0 27600 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1599_
timestamp 1644511149
transform 1 0 27784 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1600_
timestamp 1644511149
transform 1 0 29256 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1601_
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1602_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13064 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1603_
timestamp 1644511149
transform 1 0 24840 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1604_
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1605_
timestamp 1644511149
transform 1 0 29440 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1606_
timestamp 1644511149
transform 1 0 29440 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1607_
timestamp 1644511149
transform 1 0 30636 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1608_
timestamp 1644511149
transform 1 0 30820 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1609_
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1610_
timestamp 1644511149
transform 1 0 30544 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1611_
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1612_
timestamp 1644511149
transform 1 0 30820 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1613_
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1614_
timestamp 1644511149
transform 1 0 21528 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1615_
timestamp 1644511149
transform 1 0 27048 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1616_
timestamp 1644511149
transform 1 0 26312 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1617_
timestamp 1644511149
transform 1 0 26128 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1618_
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_1  _1619_
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1620_
timestamp 1644511149
transform 1 0 26036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1621_
timestamp 1644511149
transform 1 0 20976 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1622_
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1623_
timestamp 1644511149
transform 1 0 22172 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1624_
timestamp 1644511149
transform 1 0 22816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1625_
timestamp 1644511149
transform 1 0 9108 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1626_
timestamp 1644511149
transform 1 0 17020 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_1  _1627_
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1628_
timestamp 1644511149
transform 1 0 15456 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1629_
timestamp 1644511149
transform 1 0 18492 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1630_
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1631_
timestamp 1644511149
transform 1 0 20332 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1632_
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1633_
timestamp 1644511149
transform 1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1634_
timestamp 1644511149
transform 1 0 12696 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1635_
timestamp 1644511149
transform 1 0 10396 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1636_
timestamp 1644511149
transform 1 0 10580 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1637_
timestamp 1644511149
transform 1 0 9936 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1638_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12420 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1639_
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1640_
timestamp 1644511149
transform 1 0 11408 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1641_
timestamp 1644511149
transform 1 0 11684 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1642_
timestamp 1644511149
transform 1 0 12512 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1643_
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1644_
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1645_
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1646_
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1647_
timestamp 1644511149
transform 1 0 10580 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1648_
timestamp 1644511149
transform 1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1649_
timestamp 1644511149
transform 1 0 10396 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1650_
timestamp 1644511149
transform 1 0 9016 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1651_
timestamp 1644511149
transform 1 0 20148 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1652_
timestamp 1644511149
transform 1 0 12512 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1653_
timestamp 1644511149
transform 1 0 12512 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1654_
timestamp 1644511149
transform 1 0 12052 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1655_
timestamp 1644511149
transform 1 0 20884 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1656_
timestamp 1644511149
transform 1 0 22632 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_1  _1657_
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1658_
timestamp 1644511149
transform 1 0 13892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1659_
timestamp 1644511149
transform 1 0 14260 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1660_
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1661_
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1662_
timestamp 1644511149
transform 1 0 23552 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_1  _1663_
timestamp 1644511149
transform 1 0 15272 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1664_
timestamp 1644511149
transform 1 0 16100 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1665_
timestamp 1644511149
transform 1 0 24656 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1666_
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1667_
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1668_
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1669_
timestamp 1644511149
transform 1 0 17296 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1670_
timestamp 1644511149
transform 1 0 17204 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1671_
timestamp 1644511149
transform 1 0 19688 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1672_
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1673_
timestamp 1644511149
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1674_
timestamp 1644511149
transform 1 0 19320 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1675_
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1676_
timestamp 1644511149
transform 1 0 22172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1677_
timestamp 1644511149
transform 1 0 20700 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1678_
timestamp 1644511149
transform 1 0 20608 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1679_
timestamp 1644511149
transform 1 0 20884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1680_
timestamp 1644511149
transform 1 0 21712 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1681_
timestamp 1644511149
transform 1 0 21068 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1682_
timestamp 1644511149
transform 1 0 23920 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1683_
timestamp 1644511149
transform 1 0 23552 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1684_
timestamp 1644511149
transform 1 0 23276 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1685_
timestamp 1644511149
transform 1 0 21804 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1686_
timestamp 1644511149
transform 1 0 22264 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1687_
timestamp 1644511149
transform 1 0 25208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_1  _1688_
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1689_
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1690_
timestamp 1644511149
transform 1 0 25300 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1691_
timestamp 1644511149
transform 1 0 24472 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1692_
timestamp 1644511149
transform 1 0 25392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1693_
timestamp 1644511149
transform 1 0 24288 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_1  _1694_
timestamp 1644511149
transform 1 0 26404 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1695_
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1696_
timestamp 1644511149
transform 1 0 25852 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1697_
timestamp 1644511149
transform 1 0 27876 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1698_
timestamp 1644511149
transform 1 0 27784 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1699_
timestamp 1644511149
transform 1 0 28612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1700_
timestamp 1644511149
transform 1 0 28336 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1701_
timestamp 1644511149
transform 1 0 27876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1702_
timestamp 1644511149
transform 1 0 29624 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1703_
timestamp 1644511149
transform 1 0 29900 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1704_
timestamp 1644511149
transform 1 0 31372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1705_
timestamp 1644511149
transform 1 0 30544 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1706_
timestamp 1644511149
transform 1 0 30636 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1707_
timestamp 1644511149
transform 1 0 31832 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1708_
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1709_
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1710_
timestamp 1644511149
transform 1 0 32200 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1711_
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1712_
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1713_
timestamp 1644511149
transform 1 0 33764 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1714_
timestamp 1644511149
transform 1 0 36524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1715_
timestamp 1644511149
transform 1 0 22816 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1716_
timestamp 1644511149
transform 1 0 32936 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_1  _1717_
timestamp 1644511149
transform 1 0 33028 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1718_
timestamp 1644511149
transform 1 0 32568 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1719_
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1720_
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1721_
timestamp 1644511149
transform 1 0 34408 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1722_
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1723_
timestamp 1644511149
transform 1 0 32200 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1724_
timestamp 1644511149
transform 1 0 34592 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1725_
timestamp 1644511149
transform 1 0 34592 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1726_
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1727_
timestamp 1644511149
transform 1 0 12880 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1728_
timestamp 1644511149
transform 1 0 11592 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1729_
timestamp 1644511149
transform 1 0 12880 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1730_
timestamp 1644511149
transform 1 0 21896 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1731_
timestamp 1644511149
transform 1 0 22816 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1732_
timestamp 1644511149
transform 1 0 22448 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1733_
timestamp 1644511149
transform 1 0 13340 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1734_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12052 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1735_
timestamp 1644511149
transform 1 0 13340 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1736_
timestamp 1644511149
transform 1 0 21896 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1737_
timestamp 1644511149
transform 1 0 11684 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1738_
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1739_
timestamp 1644511149
transform 1 0 12972 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1740_
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1741_
timestamp 1644511149
transform 1 0 14720 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1742_
timestamp 1644511149
transform 1 0 14536 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1743_
timestamp 1644511149
transform 1 0 15364 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1744_
timestamp 1644511149
transform 1 0 20240 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1745_
timestamp 1644511149
transform 1 0 18308 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1746_
timestamp 1644511149
transform 1 0 17848 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1747_
timestamp 1644511149
transform 1 0 18952 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1748_
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1749_
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1750_
timestamp 1644511149
transform 1 0 20884 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1751_
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1752_
timestamp 1644511149
transform 1 0 18952 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1753_
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1754_
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1755_
timestamp 1644511149
transform 1 0 21896 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1756_
timestamp 1644511149
transform 1 0 20700 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1757_
timestamp 1644511149
transform 1 0 26864 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1758_
timestamp 1644511149
transform 1 0 21528 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1759_
timestamp 1644511149
transform 1 0 19596 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1760_
timestamp 1644511149
transform 1 0 25392 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1761_
timestamp 1644511149
transform 1 0 25300 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1762_
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1763_
timestamp 1644511149
transform 1 0 17020 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1764_
timestamp 1644511149
transform 1 0 26864 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1765_
timestamp 1644511149
transform 1 0 25392 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1766_
timestamp 1644511149
transform 1 0 27416 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1767_
timestamp 1644511149
transform 1 0 27232 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1768_
timestamp 1644511149
transform 1 0 28428 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1769_
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1770_
timestamp 1644511149
transform 1 0 27508 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1771_
timestamp 1644511149
transform 1 0 28152 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1772_
timestamp 1644511149
transform 1 0 27692 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1773_
timestamp 1644511149
transform 1 0 29532 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1774_
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1775_
timestamp 1644511149
transform 1 0 20792 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1776_
timestamp 1644511149
transform 1 0 23184 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1777_
timestamp 1644511149
transform 1 0 22632 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1778_
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1779_
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1780_
timestamp 1644511149
transform 1 0 25852 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1781_
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1782_
timestamp 1644511149
transform 1 0 28520 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1783_
timestamp 1644511149
transform 1 0 20700 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1784_
timestamp 1644511149
transform 1 0 20332 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1785_
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1786_
timestamp 1644511149
transform 1 0 20792 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1787_
timestamp 1644511149
transform 1 0 22908 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1788_
timestamp 1644511149
transform 1 0 21804 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1789_
timestamp 1644511149
transform 1 0 23184 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1790_
timestamp 1644511149
transform 1 0 23092 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1791_
timestamp 1644511149
transform 1 0 25300 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1792_
timestamp 1644511149
transform 1 0 25392 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1793_
timestamp 1644511149
transform 1 0 27784 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1794_
timestamp 1644511149
transform 1 0 27876 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1795_
timestamp 1644511149
transform 1 0 30636 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1796_
timestamp 1644511149
transform 1 0 29624 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1797_
timestamp 1644511149
transform 1 0 27692 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1798_
timestamp 1644511149
transform 1 0 27600 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1799_
timestamp 1644511149
transform 1 0 13432 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1800_
timestamp 1644511149
transform 1 0 28796 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1801_
timestamp 1644511149
transform 1 0 29716 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1802_
timestamp 1644511149
transform 1 0 25392 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1803_
timestamp 1644511149
transform 1 0 24472 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1804_
timestamp 1644511149
transform 1 0 24472 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1805_
timestamp 1644511149
transform 1 0 23644 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1806_
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1807_
timestamp 1644511149
transform 1 0 23092 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1808_
timestamp 1644511149
transform 1 0 12972 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1809_
timestamp 1644511149
transform 1 0 13064 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1810_
timestamp 1644511149
transform 1 0 12420 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1811_
timestamp 1644511149
transform 1 0 11224 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1812_
timestamp 1644511149
transform 1 0 13524 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1813_
timestamp 1644511149
transform 1 0 14076 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1814_
timestamp 1644511149
transform 1 0 20976 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1815_
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1816_
timestamp 1644511149
transform 1 0 15456 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1817_
timestamp 1644511149
transform 1 0 14904 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1818_
timestamp 1644511149
transform 1 0 12512 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1819_
timestamp 1644511149
transform 1 0 10304 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1820_
timestamp 1644511149
transform 1 0 13984 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1821_
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1822_
timestamp 1644511149
transform 1 0 15456 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1823_
timestamp 1644511149
transform 1 0 13984 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1824_
timestamp 1644511149
transform 1 0 15732 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1825_
timestamp 1644511149
transform 1 0 14904 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1826_
timestamp 1644511149
transform 1 0 10304 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1827_
timestamp 1644511149
transform 1 0 14720 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1828_
timestamp 1644511149
transform 1 0 14904 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1829_
timestamp 1644511149
transform 1 0 15548 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1830_
timestamp 1644511149
transform 1 0 11776 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1831_
timestamp 1644511149
transform 1 0 15732 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1832_
timestamp 1644511149
transform 1 0 16192 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1833_
timestamp 1644511149
transform 1 0 12696 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1834_
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1835_
timestamp 1644511149
transform 1 0 14720 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1836_
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1837_
timestamp 1644511149
transform 1 0 17664 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1838_
timestamp 1644511149
transform 1 0 17664 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1839_
timestamp 1644511149
transform 1 0 18124 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1840_
timestamp 1644511149
transform 1 0 18124 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1841_
timestamp 1644511149
transform 1 0 17664 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1842_
timestamp 1644511149
transform 1 0 20516 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1843_
timestamp 1644511149
transform 1 0 23000 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1844_
timestamp 1644511149
transform 1 0 23276 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_1  _1845_
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1846_
timestamp 1644511149
transform 1 0 19872 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1847_
timestamp 1644511149
transform 1 0 22540 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1848_
timestamp 1644511149
transform 1 0 21712 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1849_
timestamp 1644511149
transform 1 0 24748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1850_
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1851_
timestamp 1644511149
transform 1 0 23184 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1852_
timestamp 1644511149
transform 1 0 23276 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1853_
timestamp 1644511149
transform 1 0 26956 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1854_
timestamp 1644511149
transform 1 0 24564 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1855_
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1856_
timestamp 1644511149
transform 1 0 25576 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1857_
timestamp 1644511149
transform 1 0 31556 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1858_
timestamp 1644511149
transform 1 0 30452 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1859_
timestamp 1644511149
transform 1 0 30728 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1860_
timestamp 1644511149
transform 1 0 27600 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1861_
timestamp 1644511149
transform 1 0 29624 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1862_
timestamp 1644511149
transform 1 0 29716 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1863_
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1864_
timestamp 1644511149
transform 1 0 32292 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1865_
timestamp 1644511149
transform 1 0 32476 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1866_
timestamp 1644511149
transform 1 0 28612 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1867_
timestamp 1644511149
transform 1 0 33672 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1868_
timestamp 1644511149
transform 1 0 34684 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1869_
timestamp 1644511149
transform 1 0 28704 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1870_
timestamp 1644511149
transform 1 0 33580 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1871_
timestamp 1644511149
transform 1 0 33948 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1872_
timestamp 1644511149
transform 1 0 26128 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1873_
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1874_
timestamp 1644511149
transform 1 0 32200 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1875_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1876_
timestamp 1644511149
transform 1 0 12420 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1877_
timestamp 1644511149
transform 1 0 11960 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1878_
timestamp 1644511149
transform 1 0 11592 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1879_
timestamp 1644511149
transform 1 0 12788 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1880_
timestamp 1644511149
transform 1 0 12696 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1881_
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1882_
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1883_
timestamp 1644511149
transform 1 0 21160 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1884_
timestamp 1644511149
transform 1 0 14536 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1885_
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1886_
timestamp 1644511149
transform 1 0 15548 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1887_
timestamp 1644511149
transform 1 0 15456 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1888_
timestamp 1644511149
transform 1 0 15456 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1889_
timestamp 1644511149
transform 1 0 15456 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1890_
timestamp 1644511149
transform 1 0 17848 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1891_
timestamp 1644511149
transform 1 0 17296 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1892_
timestamp 1644511149
transform 1 0 20976 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1893_
timestamp 1644511149
transform 1 0 20976 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1894_
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1895_
timestamp 1644511149
transform 1 0 21896 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1896_
timestamp 1644511149
transform 1 0 22080 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1897_
timestamp 1644511149
transform 1 0 21068 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1898_
timestamp 1644511149
transform 1 0 19412 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1899_
timestamp 1644511149
transform 1 0 22632 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1900_
timestamp 1644511149
transform 1 0 23000 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1901_
timestamp 1644511149
transform 1 0 24104 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1902_
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1903_
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1904_
timestamp 1644511149
transform 1 0 26496 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1905_
timestamp 1644511149
transform 1 0 27600 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1906_
timestamp 1644511149
transform 1 0 27416 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1907_
timestamp 1644511149
transform 1 0 27048 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1908_
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1909_
timestamp 1644511149
transform 1 0 27416 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1910_
timestamp 1644511149
transform 1 0 18400 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1911_
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1912_
timestamp 1644511149
transform 1 0 28060 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1913_
timestamp 1644511149
transform 1 0 28244 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1914_
timestamp 1644511149
transform 1 0 25668 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1915_
timestamp 1644511149
transform 1 0 26496 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1916_
timestamp 1644511149
transform 1 0 25208 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1917_
timestamp 1644511149
transform 1 0 25024 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1918_
timestamp 1644511149
transform 1 0 23552 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1919_
timestamp 1644511149
transform 1 0 15916 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1920_
timestamp 1644511149
transform 1 0 17020 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1921_
timestamp 1644511149
transform 1 0 16560 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1922_
timestamp 1644511149
transform 1 0 20148 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1923_
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1924_
timestamp 1644511149
transform 1 0 18676 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1925_
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1926_
timestamp 1644511149
transform 1 0 17848 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1927_
timestamp 1644511149
transform 1 0 19596 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1928_
timestamp 1644511149
transform 1 0 20976 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1929_
timestamp 1644511149
transform 1 0 22264 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1930_
timestamp 1644511149
transform 1 0 21804 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1931_
timestamp 1644511149
transform 1 0 23092 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1932_
timestamp 1644511149
transform 1 0 23092 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1933_
timestamp 1644511149
transform 1 0 22816 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1934_
timestamp 1644511149
transform 1 0 27784 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1935_
timestamp 1644511149
transform 1 0 22540 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1936_
timestamp 1644511149
transform 1 0 28428 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1937_
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1938_
timestamp 1644511149
transform 1 0 29808 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1939_
timestamp 1644511149
transform 1 0 28980 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1940_
timestamp 1644511149
transform 1 0 30912 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1941_
timestamp 1644511149
transform 1 0 29440 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1942_
timestamp 1644511149
transform 1 0 30084 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1943_
timestamp 1644511149
transform 1 0 25944 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1944_
timestamp 1644511149
transform 1 0 26220 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1945_
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1946_
timestamp 1644511149
transform 1 0 13248 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1947_
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1948_
timestamp 1644511149
transform 1 0 14260 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1949_
timestamp 1644511149
transform 1 0 12972 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1950_
timestamp 1644511149
transform 1 0 13156 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1951_
timestamp 1644511149
transform 1 0 13340 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1952_
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1953_
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1954_
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1955_
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1956_
timestamp 1644511149
transform 1 0 13800 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1957_
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _1958_
timestamp 1644511149
transform 1 0 15180 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1959_
timestamp 1644511149
transform 1 0 10488 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__nor4_4  _1960_
timestamp 1644511149
transform 1 0 14904 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_1  _1961_
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1962_
timestamp 1644511149
transform 1 0 10764 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1963_
timestamp 1644511149
transform 1 0 9752 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1964_
timestamp 1644511149
transform 1 0 9660 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1965_
timestamp 1644511149
transform 1 0 10948 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1966_
timestamp 1644511149
transform 1 0 9844 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1967_
timestamp 1644511149
transform 1 0 10028 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1968_
timestamp 1644511149
transform 1 0 8648 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1969_
timestamp 1644511149
transform 1 0 9844 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1970_
timestamp 1644511149
transform 1 0 9384 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1971_
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1972_
timestamp 1644511149
transform 1 0 9568 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1973_
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1974_
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1975_
timestamp 1644511149
transform 1 0 14720 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1976_
timestamp 1644511149
transform 1 0 13524 0 -1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1977_
timestamp 1644511149
transform 1 0 15272 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1978_
timestamp 1644511149
transform 1 0 13156 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1979_
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1980_
timestamp 1644511149
transform 1 0 16468 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1981_
timestamp 1644511149
transform 1 0 14168 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1982_
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1983_
timestamp 1644511149
transform 1 0 14536 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1984_
timestamp 1644511149
transform 1 0 15732 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1985_
timestamp 1644511149
transform 1 0 15548 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1986_
timestamp 1644511149
transform 1 0 19596 0 1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1987_
timestamp 1644511149
transform 1 0 19412 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1988_
timestamp 1644511149
transform 1 0 19320 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1989_
timestamp 1644511149
transform 1 0 19504 0 -1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1990_
timestamp 1644511149
transform 1 0 19044 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1991_
timestamp 1644511149
transform 1 0 19872 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1992_
timestamp 1644511149
transform 1 0 20148 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1993_
timestamp 1644511149
transform 1 0 21620 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1994_
timestamp 1644511149
transform 1 0 20516 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1995_
timestamp 1644511149
transform 1 0 20884 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1996_
timestamp 1644511149
transform 1 0 21804 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1997_
timestamp 1644511149
transform 1 0 22448 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1998_
timestamp 1644511149
transform 1 0 20608 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1999_
timestamp 1644511149
transform 1 0 19688 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2000_
timestamp 1644511149
transform 1 0 19780 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2001_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2002_
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2003_
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2004_
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2005_
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2006_
timestamp 1644511149
transform 1 0 30176 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2007_
timestamp 1644511149
transform 1 0 30176 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2008_
timestamp 1644511149
transform 1 0 24380 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2009_
timestamp 1644511149
transform 1 0 12788 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2010_
timestamp 1644511149
transform 1 0 17664 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2011_
timestamp 1644511149
transform 1 0 19780 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2012_
timestamp 1644511149
transform 1 0 23092 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2013_
timestamp 1644511149
transform 1 0 25024 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2014_
timestamp 1644511149
transform 1 0 25024 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2015_
timestamp 1644511149
transform 1 0 25392 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2016_
timestamp 1644511149
transform 1 0 16836 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2017_
timestamp 1644511149
transform 1 0 9016 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2018_
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2019_
timestamp 1644511149
transform 1 0 4416 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2020_
timestamp 1644511149
transform 1 0 34500 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2021_
timestamp 1644511149
transform 1 0 3496 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2022_
timestamp 1644511149
transform 1 0 34500 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2023_
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2024_
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2025_
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2026_
timestamp 1644511149
transform 1 0 32660 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2027_
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2028_
timestamp 1644511149
transform 1 0 34684 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2029_
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2030_
timestamp 1644511149
transform 1 0 32752 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2031_
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2032_
timestamp 1644511149
transform 1 0 36524 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2033_
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2034_
timestamp 1644511149
transform 1 0 34500 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2035_
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2036_
timestamp 1644511149
transform 1 0 32660 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2037_
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2038_
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2039_
timestamp 1644511149
transform 1 0 5612 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2040_
timestamp 1644511149
transform 1 0 32660 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2041_
timestamp 1644511149
transform 1 0 6164 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2042_
timestamp 1644511149
transform 1 0 32660 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2043_
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2044_
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2045_
timestamp 1644511149
transform 1 0 8188 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2046_
timestamp 1644511149
transform 1 0 32660 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2047_
timestamp 1644511149
transform 1 0 3864 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2048_
timestamp 1644511149
transform 1 0 29900 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2049_
timestamp 1644511149
transform 1 0 6992 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2050_
timestamp 1644511149
transform 1 0 2668 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2051_
timestamp 1644511149
transform 1 0 7176 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2052_
timestamp 1644511149
transform 1 0 2668 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2053_
timestamp 1644511149
transform 1 0 4968 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2054_
timestamp 1644511149
transform 1 0 1840 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2055_
timestamp 1644511149
transform 1 0 4968 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2056_
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2057_
timestamp 1644511149
transform 1 0 5336 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2058_
timestamp 1644511149
transform 1 0 7360 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2059_
timestamp 1644511149
transform 1 0 7268 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2060_
timestamp 1644511149
transform 1 0 2668 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2061_
timestamp 1644511149
transform 1 0 9108 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2062_
timestamp 1644511149
transform 1 0 2668 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2063_
timestamp 1644511149
transform 1 0 6992 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2064_
timestamp 1644511149
transform 1 0 1840 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2065_
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2066_
timestamp 1644511149
transform 1 0 1840 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2067_
timestamp 1644511149
transform 1 0 4416 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2068_
timestamp 1644511149
transform 1 0 6992 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2069_
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2070_
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2071_
timestamp 1644511149
transform 1 0 8924 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2072_
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2073_
timestamp 1644511149
transform 1 0 9292 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2074_
timestamp 1644511149
transform 1 0 5612 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2075_
timestamp 1644511149
transform 1 0 10764 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2076_
timestamp 1644511149
transform 1 0 2668 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2077_
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2078_
timestamp 1644511149
transform 1 0 6992 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2079_
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2080_
timestamp 1644511149
transform 1 0 7912 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2081_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2082_
timestamp 1644511149
transform 1 0 7912 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2083_
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2084_
timestamp 1644511149
transform 1 0 6808 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2085_
timestamp 1644511149
transform 1 0 8648 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2086_
timestamp 1644511149
transform 1 0 9752 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2087_
timestamp 1644511149
transform 1 0 9752 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2088_
timestamp 1644511149
transform 1 0 11684 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2089_
timestamp 1644511149
transform 1 0 12052 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2090_
timestamp 1644511149
transform 1 0 14628 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2091_
timestamp 1644511149
transform 1 0 12052 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2092_
timestamp 1644511149
transform 1 0 17204 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2093_
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2094_
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2095_
timestamp 1644511149
transform 1 0 20424 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2096_
timestamp 1644511149
transform 1 0 20516 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2097_
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2098_
timestamp 1644511149
transform 1 0 21896 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2099_
timestamp 1644511149
transform 1 0 23736 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2100_
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2101_
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2102_
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2103_
timestamp 1644511149
transform 1 0 27140 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2104_
timestamp 1644511149
transform 1 0 27508 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2105_
timestamp 1644511149
transform 1 0 28520 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2106_
timestamp 1644511149
transform 1 0 29900 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2107_
timestamp 1644511149
transform 1 0 29992 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2108_
timestamp 1644511149
transform 1 0 30084 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2109_
timestamp 1644511149
transform 1 0 31004 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2110_
timestamp 1644511149
transform 1 0 25024 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2111_
timestamp 1644511149
transform 1 0 25576 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2112_
timestamp 1644511149
transform 1 0 22356 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2113_
timestamp 1644511149
transform 1 0 16100 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2114_
timestamp 1644511149
transform 1 0 20240 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2115_
timestamp 1644511149
transform 1 0 8372 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2116_
timestamp 1644511149
transform 1 0 9844 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2117_
timestamp 1644511149
transform 1 0 13524 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2118_
timestamp 1644511149
transform 1 0 11684 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2119_
timestamp 1644511149
transform 1 0 7544 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2120_
timestamp 1644511149
transform 1 0 9752 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2121_
timestamp 1644511149
transform 1 0 8556 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2122_
timestamp 1644511149
transform 1 0 11592 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2123_
timestamp 1644511149
transform 1 0 12512 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2124_
timestamp 1644511149
transform 1 0 13432 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2125_
timestamp 1644511149
transform 1 0 14628 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2126_
timestamp 1644511149
transform 1 0 15456 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2127_
timestamp 1644511149
transform 1 0 16836 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2128_
timestamp 1644511149
transform 1 0 17848 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2129_
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2130_
timestamp 1644511149
transform 1 0 19964 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2131_
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2132_
timestamp 1644511149
transform 1 0 22448 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2133_
timestamp 1644511149
transform 1 0 23368 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2134_
timestamp 1644511149
transform 1 0 25024 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2135_
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2136_
timestamp 1644511149
transform 1 0 27324 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2137_
timestamp 1644511149
transform 1 0 28796 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2138_
timestamp 1644511149
transform 1 0 29624 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2139_
timestamp 1644511149
transform 1 0 30084 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2140_
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2141_
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2142_
timestamp 1644511149
transform 1 0 33948 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2143_
timestamp 1644511149
transform 1 0 32384 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2144_
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2145_
timestamp 1644511149
transform 1 0 32568 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2146_
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2147_
timestamp 1644511149
transform 1 0 12696 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2148_
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2149_
timestamp 1644511149
transform 1 0 14628 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2150_
timestamp 1644511149
transform 1 0 12144 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2151_
timestamp 1644511149
transform 1 0 15364 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2152_
timestamp 1644511149
transform 1 0 18400 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2153_
timestamp 1644511149
transform 1 0 18584 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2154_
timestamp 1644511149
transform 1 0 22172 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2155_
timestamp 1644511149
transform 1 0 21896 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2156_
timestamp 1644511149
transform 1 0 24932 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2157_
timestamp 1644511149
transform 1 0 25024 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2158_
timestamp 1644511149
transform 1 0 27508 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2159_
timestamp 1644511149
transform 1 0 29808 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2160_
timestamp 1644511149
transform 1 0 27600 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2161_
timestamp 1644511149
transform 1 0 29992 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2162_
timestamp 1644511149
transform 1 0 20608 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2163_
timestamp 1644511149
transform 1 0 22448 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2164_
timestamp 1644511149
transform 1 0 17296 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2165_
timestamp 1644511149
transform 1 0 19228 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2166_
timestamp 1644511149
transform 1 0 20608 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2167_
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2168_
timestamp 1644511149
transform 1 0 22448 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2169_
timestamp 1644511149
transform 1 0 25392 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2170_
timestamp 1644511149
transform 1 0 28888 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2171_
timestamp 1644511149
transform 1 0 30084 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2172_
timestamp 1644511149
transform 1 0 27508 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2173_
timestamp 1644511149
transform 1 0 31924 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2174_
timestamp 1644511149
transform 1 0 24932 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2175_
timestamp 1644511149
transform 1 0 23184 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2176_
timestamp 1644511149
transform 1 0 11224 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2177_
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2178_
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2179_
timestamp 1644511149
transform 1 0 14628 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2180_
timestamp 1644511149
transform 1 0 10948 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2181_
timestamp 1644511149
transform 1 0 14260 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2182_
timestamp 1644511149
transform 1 0 9752 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2183_
timestamp 1644511149
transform 1 0 14628 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2184_
timestamp 1644511149
transform 1 0 9568 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2185_
timestamp 1644511149
transform 1 0 16468 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2186_
timestamp 1644511149
transform 1 0 12144 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2187_
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2188_
timestamp 1644511149
transform 1 0 14076 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2189_
timestamp 1644511149
transform 1 0 16744 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2190_
timestamp 1644511149
transform 1 0 17296 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2191_
timestamp 1644511149
transform 1 0 17388 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2192_
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2193_
timestamp 1644511149
transform 1 0 21160 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2194_
timestamp 1644511149
transform 1 0 19872 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2195_
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2196_
timestamp 1644511149
transform 1 0 22816 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2197_
timestamp 1644511149
transform 1 0 22448 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2198_
timestamp 1644511149
transform 1 0 24748 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2199_
timestamp 1644511149
transform 1 0 24840 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2200_
timestamp 1644511149
transform 1 0 25576 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2201_
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2202_
timestamp 1644511149
transform 1 0 27232 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2203_
timestamp 1644511149
transform 1 0 29716 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2204_
timestamp 1644511149
transform 1 0 27140 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2205_
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2206_
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2207_
timestamp 1644511149
transform 1 0 33764 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2208_
timestamp 1644511149
transform 1 0 27876 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2209_
timestamp 1644511149
transform 1 0 33580 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2210_
timestamp 1644511149
transform 1 0 25024 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2211_
timestamp 1644511149
transform 1 0 32292 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2212_
timestamp 1644511149
transform 1 0 19044 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2213_
timestamp 1644511149
transform 1 0 12052 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2214_
timestamp 1644511149
transform 1 0 10120 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2215_
timestamp 1644511149
transform 1 0 12696 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2216_
timestamp 1644511149
transform 1 0 14536 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2217_
timestamp 1644511149
transform 1 0 15732 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2218_
timestamp 1644511149
transform 1 0 16008 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2219_
timestamp 1644511149
transform 1 0 17480 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2220_
timestamp 1644511149
transform 1 0 21896 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2221_
timestamp 1644511149
transform 1 0 22356 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2222_
timestamp 1644511149
transform 1 0 22264 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2223_
timestamp 1644511149
transform 1 0 24104 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2224_
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2225_
timestamp 1644511149
transform 1 0 28796 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2226_
timestamp 1644511149
transform 1 0 27416 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2227_
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2228_
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2229_
timestamp 1644511149
transform 1 0 25024 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2230_
timestamp 1644511149
transform 1 0 17388 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2231_
timestamp 1644511149
transform 1 0 16836 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2232_
timestamp 1644511149
transform 1 0 19228 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2233_
timestamp 1644511149
transform 1 0 19688 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2234_
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2235_
timestamp 1644511149
transform 1 0 22448 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2236_
timestamp 1644511149
transform 1 0 29532 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2237_
timestamp 1644511149
transform 1 0 30544 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2238_
timestamp 1644511149
transform 1 0 30176 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2239_
timestamp 1644511149
transform 1 0 31372 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2240_
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2241_
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2242_
timestamp 1644511149
transform 1 0 12972 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2243_
timestamp 1644511149
transform 1 0 14076 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2244_
timestamp 1644511149
transform 1 0 14260 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2245_
timestamp 1644511149
transform 1 0 15456 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2246_
timestamp 1644511149
transform 1 0 9568 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2247_
timestamp 1644511149
transform 1 0 9568 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2248_
timestamp 1644511149
transform 1 0 9292 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2249_
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2250_
timestamp 1644511149
transform 1 0 9200 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2251_
timestamp 1644511149
transform 1 0 15640 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2252_
timestamp 1644511149
transform 1 0 12696 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2253_
timestamp 1644511149
transform 1 0 14720 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2254_
timestamp 1644511149
transform 1 0 12880 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2255_
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2256_
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2257_
timestamp 1644511149
transform 1 0 19780 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2258_
timestamp 1644511149
transform 1 0 20884 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2259_
timestamp 1644511149
transform 1 0 21896 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2260_
timestamp 1644511149
transform 1 0 21988 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2261_
timestamp 1644511149
transform 1 0 19780 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _2262__150 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2263__151
timestamp 1644511149
transform 1 0 2116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CLK pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19412 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_CLK
timestamp 1644511149
transform 1 0 19872 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_CLK
timestamp 1644511149
transform 1 0 18032 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_CLK
timestamp 1644511149
transform 1 0 9200 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_CLK
timestamp 1644511149
transform 1 0 28980 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_CLK
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_CLK
timestamp 1644511149
transform 1 0 29348 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_CLK
timestamp 1644511149
transform 1 0 5612 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_CLK
timestamp 1644511149
transform 1 0 4140 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_CLK
timestamp 1644511149
transform 1 0 9200 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_CLK
timestamp 1644511149
transform 1 0 11868 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_CLK
timestamp 1644511149
transform 1 0 15548 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_CLK
timestamp 1644511149
transform 1 0 10488 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_CLK
timestamp 1644511149
transform 1 0 5520 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_CLK
timestamp 1644511149
transform 1 0 10672 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_CLK
timestamp 1644511149
transform 1 0 15824 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_CLK
timestamp 1644511149
transform 1 0 15640 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_CLK
timestamp 1644511149
transform 1 0 20608 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_11_CLK
timestamp 1644511149
transform 1 0 25668 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_12_CLK
timestamp 1644511149
transform 1 0 21252 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_13_CLK
timestamp 1644511149
transform 1 0 27232 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_14_CLK
timestamp 1644511149
transform 1 0 31096 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_15_CLK
timestamp 1644511149
transform 1 0 27324 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_16_CLK
timestamp 1644511149
transform 1 0 24012 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_17_CLK
timestamp 1644511149
transform 1 0 30084 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_18_CLK
timestamp 1644511149
transform 1 0 35052 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_19_CLK
timestamp 1644511149
transform 1 0 32384 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_20_CLK
timestamp 1644511149
transform 1 0 32292 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_21_CLK
timestamp 1644511149
transform 1 0 26404 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_22_CLK
timestamp 1644511149
transform 1 0 22172 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_23_CLK
timestamp 1644511149
transform 1 0 24748 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_24_CLK
timestamp 1644511149
transform 1 0 19136 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_25_CLK
timestamp 1644511149
transform 1 0 14352 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_26_CLK
timestamp 1644511149
transform 1 0 14352 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_27_CLK
timestamp 1644511149
transform 1 0 9200 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17756 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1644511149
transform 1 0 21896 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19872 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1644511149
transform 1 0 1656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1644511149
transform 1 0 27324 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1644511149
transform 1 0 35144 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1644511149
transform 1 0 35880 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1644511149
transform 1 0 37076 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1644511149
transform 1 0 37260 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1644511149
transform 1 0 37812 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1644511149
transform 1 0 28060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1644511149
transform 1 0 29624 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1644511149
transform 1 0 32108 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1644511149
transform 1 0 31280 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1644511149
transform 1 0 32936 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1644511149
transform 1 0 33764 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1644511149
transform 1 0 34592 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1644511149
transform 1 0 3772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1644511149
transform 1 0 17296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1644511149
transform 1 0 18124 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform 1 0 18032 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform 1 0 19872 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform 1 0 20240 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1644511149
transform 1 0 22908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1644511149
transform 1 0 23552 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 27232 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 28428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform 1 0 4600 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform 1 0 27140 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1644511149
transform 1 0 32752 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1644511149
transform 1 0 33396 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1644511149
transform 1 0 33580 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1644511149
transform 1 0 35144 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1644511149
transform 1 0 35788 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1644511149
transform 1 0 37168 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1644511149
transform 1 0 37904 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1644511149
transform 1 0 7636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1644511149
transform 1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1644511149
transform 1 0 10212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1644511149
transform 1 0 11316 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1644511149
transform 1 0 12696 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1644511149
transform 1 0 16468 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1644511149
transform 1 0 17112 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1644511149
transform 1 0 17756 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1644511149
transform 1 0 17480 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1644511149
transform 1 0 18676 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1644511149
transform 1 0 19504 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1644511149
transform 1 0 25024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1644511149
transform 1 0 25668 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1644511149
transform 1 0 28612 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1644511149
transform 1 0 4968 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1644511149
transform 1 0 30176 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1644511149
transform 1 0 30912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1644511149
transform 1 0 30820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1644511149
transform 1 0 31464 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1644511149
transform 1 0 31556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1644511149
transform 1 0 33856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1644511149
transform 1 0 35696 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1644511149
transform 1 0 35052 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input71
timestamp 1644511149
transform 1 0 35880 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input72
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1644511149
transform 1 0 6532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1644511149
transform 1 0 37812 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1644511149
transform 1 0 7544 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1644511149
transform 1 0 9476 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1644511149
transform 1 0 10580 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1644511149
transform 1 0 11684 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1644511149
transform 1 0 13524 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1644511149
transform 1 0 14168 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1644511149
transform 1 0 15088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1644511149
transform 1 0 2484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input84
timestamp 1644511149
transform 1 0 2392 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1644511149
transform 1 0 9660 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1644511149
transform 1 0 10396 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1644511149
transform 1 0 11500 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1644511149
transform 1 0 12236 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1644511149
transform 1 0 12972 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1644511149
transform 1 0 2116 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1644511149
transform 1 0 2852 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1644511149
transform 1 0 4508 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1644511149
transform 1 0 5244 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1644511149
transform 1 0 5428 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1644511149
transform 1 0 6348 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1644511149
transform 1 0 7084 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1644511149
transform 1 0 7912 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1644511149
transform 1 0 22080 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1644511149
transform 1 0 22908 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1644511149
transform 1 0 25116 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1644511149
transform 1 0 25852 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1644511149
transform 1 0 14812 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1644511149
transform 1 0 15548 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1644511149
transform 1 0 16652 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1644511149
transform 1 0 17388 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1644511149
transform 1 0 18124 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1644511149
transform 1 0 19964 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1644511149
transform 1 0 20700 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1644511149
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1644511149
transform 1 0 15824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1644511149
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1644511149
transform 1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1644511149
transform 1 0 22540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1644511149
transform 1 0 23276 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1644511149
transform 1 0 25944 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1644511149
transform 1 0 5428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1644511149
transform 1 0 27692 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1644511149
transform 1 0 30728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1644511149
transform 1 0 32936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1644511149
transform 1 0 33672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1644511149
transform 1 0 35788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1644511149
transform 1 0 35696 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1644511149
transform 1 0 36524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1644511149
transform 1 0 37628 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1644511149
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1644511149
transform 1 0 37812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1644511149
transform 1 0 37812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1644511149
transform 1 0 9844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1644511149
transform 1 0 12236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1644511149
transform 1 0 13156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1644511149
transform 1 0 15272 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1644511149
transform 1 0 14628 0 -1 4352
box -38 -48 406 592
<< labels >>
rlabel metal2 s 202 0 258 800 6 CLK
port 0 nsew signal input
rlabel metal2 s 570 0 626 800 6 RST_N
port 1 nsew signal input
rlabel metal2 s 27066 49200 27122 50000 6 in[0]
port 2 nsew signal input
rlabel metal2 s 35346 49200 35402 50000 6 in[10]
port 3 nsew signal input
rlabel metal2 s 36174 49200 36230 50000 6 in[11]
port 4 nsew signal input
rlabel metal2 s 37002 49200 37058 50000 6 in[12]
port 5 nsew signal input
rlabel metal2 s 37830 49200 37886 50000 6 in[13]
port 6 nsew signal input
rlabel metal2 s 38658 49200 38714 50000 6 in[14]
port 7 nsew signal input
rlabel metal2 s 39486 49200 39542 50000 6 in[15]
port 8 nsew signal input
rlabel metal2 s 27894 49200 27950 50000 6 in[1]
port 9 nsew signal input
rlabel metal2 s 28722 49200 28778 50000 6 in[2]
port 10 nsew signal input
rlabel metal2 s 29550 49200 29606 50000 6 in[3]
port 11 nsew signal input
rlabel metal2 s 30378 49200 30434 50000 6 in[4]
port 12 nsew signal input
rlabel metal2 s 31206 49200 31262 50000 6 in[5]
port 13 nsew signal input
rlabel metal2 s 32034 49200 32090 50000 6 in[6]
port 14 nsew signal input
rlabel metal2 s 32862 49200 32918 50000 6 in[7]
port 15 nsew signal input
rlabel metal2 s 33690 49200 33746 50000 6 in[8]
port 16 nsew signal input
rlabel metal2 s 34518 49200 34574 50000 6 in[9]
port 17 nsew signal input
rlabel metal2 s 386 49200 442 50000 6 oe[0]
port 18 nsew signal tristate
rlabel metal2 s 8666 49200 8722 50000 6 oe[10]
port 19 nsew signal tristate
rlabel metal2 s 9494 49200 9550 50000 6 oe[11]
port 20 nsew signal tristate
rlabel metal2 s 10322 49200 10378 50000 6 oe[12]
port 21 nsew signal tristate
rlabel metal2 s 11150 49200 11206 50000 6 oe[13]
port 22 nsew signal tristate
rlabel metal2 s 11978 49200 12034 50000 6 oe[14]
port 23 nsew signal tristate
rlabel metal2 s 12806 49200 12862 50000 6 oe[15]
port 24 nsew signal tristate
rlabel metal2 s 1214 49200 1270 50000 6 oe[1]
port 25 nsew signal tristate
rlabel metal2 s 2042 49200 2098 50000 6 oe[2]
port 26 nsew signal tristate
rlabel metal2 s 2870 49200 2926 50000 6 oe[3]
port 27 nsew signal tristate
rlabel metal2 s 3698 49200 3754 50000 6 oe[4]
port 28 nsew signal tristate
rlabel metal2 s 4526 49200 4582 50000 6 oe[5]
port 29 nsew signal tristate
rlabel metal2 s 5354 49200 5410 50000 6 oe[6]
port 30 nsew signal tristate
rlabel metal2 s 6182 49200 6238 50000 6 oe[7]
port 31 nsew signal tristate
rlabel metal2 s 7010 49200 7066 50000 6 oe[8]
port 32 nsew signal tristate
rlabel metal2 s 7838 49200 7894 50000 6 oe[9]
port 33 nsew signal tristate
rlabel metal2 s 13726 49200 13782 50000 6 out[0]
port 34 nsew signal tristate
rlabel metal2 s 22006 49200 22062 50000 6 out[10]
port 35 nsew signal tristate
rlabel metal2 s 22834 49200 22890 50000 6 out[11]
port 36 nsew signal tristate
rlabel metal2 s 23662 49200 23718 50000 6 out[12]
port 37 nsew signal tristate
rlabel metal2 s 24490 49200 24546 50000 6 out[13]
port 38 nsew signal tristate
rlabel metal2 s 25318 49200 25374 50000 6 out[14]
port 39 nsew signal tristate
rlabel metal2 s 26146 49200 26202 50000 6 out[15]
port 40 nsew signal tristate
rlabel metal2 s 14554 49200 14610 50000 6 out[1]
port 41 nsew signal tristate
rlabel metal2 s 15382 49200 15438 50000 6 out[2]
port 42 nsew signal tristate
rlabel metal2 s 16210 49200 16266 50000 6 out[3]
port 43 nsew signal tristate
rlabel metal2 s 17038 49200 17094 50000 6 out[4]
port 44 nsew signal tristate
rlabel metal2 s 17866 49200 17922 50000 6 out[5]
port 45 nsew signal tristate
rlabel metal2 s 18694 49200 18750 50000 6 out[6]
port 46 nsew signal tristate
rlabel metal2 s 19522 49200 19578 50000 6 out[7]
port 47 nsew signal tristate
rlabel metal2 s 20350 49200 20406 50000 6 out[8]
port 48 nsew signal tristate
rlabel metal2 s 21178 49200 21234 50000 6 out[9]
port 49 nsew signal tristate
rlabel metal2 s 938 0 994 800 6 slave_ack_o
port 50 nsew signal tristate
rlabel metal2 s 3146 0 3202 800 6 slave_adr_i[0]
port 51 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 slave_adr_i[10]
port 52 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 slave_adr_i[11]
port 53 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 slave_adr_i[12]
port 54 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 slave_adr_i[13]
port 55 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 slave_adr_i[14]
port 56 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 slave_adr_i[15]
port 57 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 slave_adr_i[16]
port 58 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 slave_adr_i[17]
port 59 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 slave_adr_i[18]
port 60 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 slave_adr_i[19]
port 61 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 slave_adr_i[1]
port 62 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 slave_adr_i[20]
port 63 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 slave_adr_i[21]
port 64 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 slave_adr_i[22]
port 65 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 slave_adr_i[23]
port 66 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 slave_adr_i[24]
port 67 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 slave_adr_i[25]
port 68 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 slave_adr_i[26]
port 69 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 slave_adr_i[27]
port 70 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 slave_adr_i[28]
port 71 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 slave_adr_i[29]
port 72 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 slave_adr_i[2]
port 73 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 slave_adr_i[30]
port 74 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 slave_adr_i[31]
port 75 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 slave_adr_i[3]
port 76 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 slave_adr_i[4]
port 77 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 slave_adr_i[5]
port 78 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 slave_adr_i[6]
port 79 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 slave_adr_i[7]
port 80 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 slave_adr_i[8]
port 81 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 slave_adr_i[9]
port 82 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 slave_cyc_i
port 83 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 slave_dat_i[0]
port 84 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 slave_dat_i[10]
port 85 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 slave_dat_i[11]
port 86 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 slave_dat_i[12]
port 87 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 slave_dat_i[13]
port 88 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 slave_dat_i[14]
port 89 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 slave_dat_i[15]
port 90 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 slave_dat_i[16]
port 91 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 slave_dat_i[17]
port 92 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 slave_dat_i[18]
port 93 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 slave_dat_i[19]
port 94 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 slave_dat_i[1]
port 95 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 slave_dat_i[20]
port 96 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 slave_dat_i[21]
port 97 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 slave_dat_i[22]
port 98 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 slave_dat_i[23]
port 99 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 slave_dat_i[24]
port 100 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 slave_dat_i[25]
port 101 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 slave_dat_i[26]
port 102 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 slave_dat_i[27]
port 103 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 slave_dat_i[28]
port 104 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 slave_dat_i[29]
port 105 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 slave_dat_i[2]
port 106 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 slave_dat_i[30]
port 107 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 slave_dat_i[31]
port 108 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 slave_dat_i[3]
port 109 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 slave_dat_i[4]
port 110 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 slave_dat_i[5]
port 111 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 slave_dat_i[6]
port 112 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 slave_dat_i[7]
port 113 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 slave_dat_i[8]
port 114 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 slave_dat_i[9]
port 115 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 slave_dat_o[0]
port 116 nsew signal tristate
rlabel metal2 s 16486 0 16542 800 6 slave_dat_o[10]
port 117 nsew signal tristate
rlabel metal2 s 17590 0 17646 800 6 slave_dat_o[11]
port 118 nsew signal tristate
rlabel metal2 s 18694 0 18750 800 6 slave_dat_o[12]
port 119 nsew signal tristate
rlabel metal2 s 19798 0 19854 800 6 slave_dat_o[13]
port 120 nsew signal tristate
rlabel metal2 s 20902 0 20958 800 6 slave_dat_o[14]
port 121 nsew signal tristate
rlabel metal2 s 22006 0 22062 800 6 slave_dat_o[15]
port 122 nsew signal tristate
rlabel metal2 s 23110 0 23166 800 6 slave_dat_o[16]
port 123 nsew signal tristate
rlabel metal2 s 24214 0 24270 800 6 slave_dat_o[17]
port 124 nsew signal tristate
rlabel metal2 s 25318 0 25374 800 6 slave_dat_o[18]
port 125 nsew signal tristate
rlabel metal2 s 26422 0 26478 800 6 slave_dat_o[19]
port 126 nsew signal tristate
rlabel metal2 s 5354 0 5410 800 6 slave_dat_o[1]
port 127 nsew signal tristate
rlabel metal2 s 27618 0 27674 800 6 slave_dat_o[20]
port 128 nsew signal tristate
rlabel metal2 s 28722 0 28778 800 6 slave_dat_o[21]
port 129 nsew signal tristate
rlabel metal2 s 29826 0 29882 800 6 slave_dat_o[22]
port 130 nsew signal tristate
rlabel metal2 s 30930 0 30986 800 6 slave_dat_o[23]
port 131 nsew signal tristate
rlabel metal2 s 32034 0 32090 800 6 slave_dat_o[24]
port 132 nsew signal tristate
rlabel metal2 s 33138 0 33194 800 6 slave_dat_o[25]
port 133 nsew signal tristate
rlabel metal2 s 34242 0 34298 800 6 slave_dat_o[26]
port 134 nsew signal tristate
rlabel metal2 s 35346 0 35402 800 6 slave_dat_o[27]
port 135 nsew signal tristate
rlabel metal2 s 36450 0 36506 800 6 slave_dat_o[28]
port 136 nsew signal tristate
rlabel metal2 s 37554 0 37610 800 6 slave_dat_o[29]
port 137 nsew signal tristate
rlabel metal2 s 6826 0 6882 800 6 slave_dat_o[2]
port 138 nsew signal tristate
rlabel metal2 s 38658 0 38714 800 6 slave_dat_o[30]
port 139 nsew signal tristate
rlabel metal2 s 39762 0 39818 800 6 slave_dat_o[31]
port 140 nsew signal tristate
rlabel metal2 s 8298 0 8354 800 6 slave_dat_o[3]
port 141 nsew signal tristate
rlabel metal2 s 9770 0 9826 800 6 slave_dat_o[4]
port 142 nsew signal tristate
rlabel metal2 s 10874 0 10930 800 6 slave_dat_o[5]
port 143 nsew signal tristate
rlabel metal2 s 11978 0 12034 800 6 slave_dat_o[6]
port 144 nsew signal tristate
rlabel metal2 s 13082 0 13138 800 6 slave_dat_o[7]
port 145 nsew signal tristate
rlabel metal2 s 14278 0 14334 800 6 slave_dat_o[8]
port 146 nsew signal tristate
rlabel metal2 s 15382 0 15438 800 6 slave_dat_o[9]
port 147 nsew signal tristate
rlabel metal2 s 1674 0 1730 800 6 slave_err_o
port 148 nsew signal tristate
rlabel metal2 s 2042 0 2098 800 6 slave_rty_o
port 149 nsew signal tristate
rlabel metal2 s 4250 0 4306 800 6 slave_sel_i[0]
port 150 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 slave_sel_i[1]
port 151 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 slave_sel_i[2]
port 152 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 slave_sel_i[3]
port 153 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 slave_stb_i
port 154 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 slave_we_i
port 155 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 156 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 156 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 157 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 40000 50000
<< end >>
