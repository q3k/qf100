VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mkQF100Fabric
  CLASS BLOCK ;
  FOREIGN mkQF100Fabric ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 300.000 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END CLK
  PIN RST_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END RST_N
  PIN cpu_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END cpu_ack_o
  PIN cpu_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END cpu_adr_i[0]
  PIN cpu_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END cpu_adr_i[10]
  PIN cpu_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END cpu_adr_i[11]
  PIN cpu_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END cpu_adr_i[12]
  PIN cpu_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END cpu_adr_i[13]
  PIN cpu_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END cpu_adr_i[14]
  PIN cpu_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END cpu_adr_i[15]
  PIN cpu_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END cpu_adr_i[16]
  PIN cpu_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.160 4.000 176.760 ;
    END
  END cpu_adr_i[17]
  PIN cpu_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END cpu_adr_i[18]
  PIN cpu_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END cpu_adr_i[19]
  PIN cpu_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END cpu_adr_i[1]
  PIN cpu_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END cpu_adr_i[20]
  PIN cpu_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END cpu_adr_i[21]
  PIN cpu_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END cpu_adr_i[22]
  PIN cpu_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END cpu_adr_i[23]
  PIN cpu_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END cpu_adr_i[24]
  PIN cpu_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.800 4.000 243.400 ;
    END
  END cpu_adr_i[25]
  PIN cpu_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.960 4.000 251.560 ;
    END
  END cpu_adr_i[26]
  PIN cpu_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END cpu_adr_i[27]
  PIN cpu_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END cpu_adr_i[28]
  PIN cpu_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END cpu_adr_i[29]
  PIN cpu_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END cpu_adr_i[2]
  PIN cpu_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END cpu_adr_i[30]
  PIN cpu_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END cpu_adr_i[31]
  PIN cpu_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END cpu_adr_i[3]
  PIN cpu_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END cpu_adr_i[4]
  PIN cpu_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END cpu_adr_i[5]
  PIN cpu_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END cpu_adr_i[6]
  PIN cpu_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END cpu_adr_i[7]
  PIN cpu_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END cpu_adr_i[8]
  PIN cpu_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END cpu_adr_i[9]
  PIN cpu_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END cpu_cyc_i
  PIN cpu_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END cpu_dat_i[0]
  PIN cpu_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END cpu_dat_i[10]
  PIN cpu_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 4.000 129.160 ;
    END
  END cpu_dat_i[11]
  PIN cpu_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END cpu_dat_i[12]
  PIN cpu_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END cpu_dat_i[13]
  PIN cpu_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END cpu_dat_i[14]
  PIN cpu_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END cpu_dat_i[15]
  PIN cpu_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END cpu_dat_i[16]
  PIN cpu_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END cpu_dat_i[17]
  PIN cpu_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END cpu_dat_i[18]
  PIN cpu_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END cpu_dat_i[19]
  PIN cpu_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END cpu_dat_i[1]
  PIN cpu_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END cpu_dat_i[20]
  PIN cpu_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END cpu_dat_i[21]
  PIN cpu_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END cpu_dat_i[22]
  PIN cpu_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END cpu_dat_i[23]
  PIN cpu_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.360 4.000 237.960 ;
    END
  END cpu_dat_i[24]
  PIN cpu_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END cpu_dat_i[25]
  PIN cpu_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.680 4.000 254.280 ;
    END
  END cpu_dat_i[26]
  PIN cpu_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END cpu_dat_i[27]
  PIN cpu_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END cpu_dat_i[28]
  PIN cpu_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END cpu_dat_i[29]
  PIN cpu_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END cpu_dat_i[2]
  PIN cpu_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END cpu_dat_i[30]
  PIN cpu_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END cpu_dat_i[31]
  PIN cpu_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END cpu_dat_i[3]
  PIN cpu_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END cpu_dat_i[4]
  PIN cpu_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END cpu_dat_i[5]
  PIN cpu_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END cpu_dat_i[6]
  PIN cpu_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END cpu_dat_i[7]
  PIN cpu_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 4.000 104.680 ;
    END
  END cpu_dat_i[8]
  PIN cpu_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END cpu_dat_i[9]
  PIN cpu_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END cpu_dat_o[0]
  PIN cpu_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END cpu_dat_o[10]
  PIN cpu_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END cpu_dat_o[11]
  PIN cpu_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END cpu_dat_o[12]
  PIN cpu_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END cpu_dat_o[13]
  PIN cpu_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END cpu_dat_o[14]
  PIN cpu_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END cpu_dat_o[15]
  PIN cpu_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END cpu_dat_o[16]
  PIN cpu_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.600 4.000 182.200 ;
    END
  END cpu_dat_o[17]
  PIN cpu_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.760 4.000 190.360 ;
    END
  END cpu_dat_o[18]
  PIN cpu_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END cpu_dat_o[19]
  PIN cpu_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END cpu_dat_o[1]
  PIN cpu_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END cpu_dat_o[20]
  PIN cpu_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END cpu_dat_o[21]
  PIN cpu_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END cpu_dat_o[22]
  PIN cpu_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END cpu_dat_o[23]
  PIN cpu_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END cpu_dat_o[24]
  PIN cpu_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END cpu_dat_o[25]
  PIN cpu_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.400 4.000 257.000 ;
    END
  END cpu_dat_o[26]
  PIN cpu_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END cpu_dat_o[27]
  PIN cpu_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END cpu_dat_o[28]
  PIN cpu_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END cpu_dat_o[29]
  PIN cpu_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END cpu_dat_o[2]
  PIN cpu_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END cpu_dat_o[30]
  PIN cpu_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END cpu_dat_o[31]
  PIN cpu_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END cpu_dat_o[3]
  PIN cpu_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END cpu_dat_o[4]
  PIN cpu_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END cpu_dat_o[5]
  PIN cpu_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END cpu_dat_o[6]
  PIN cpu_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END cpu_dat_o[7]
  PIN cpu_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END cpu_dat_o[8]
  PIN cpu_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END cpu_dat_o[9]
  PIN cpu_err_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END cpu_err_o
  PIN cpu_rty_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END cpu_rty_o
  PIN cpu_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END cpu_sel_i[0]
  PIN cpu_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END cpu_sel_i[1]
  PIN cpu_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END cpu_sel_i[2]
  PIN cpu_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END cpu_sel_i[3]
  PIN cpu_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END cpu_stb_i
  PIN cpu_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END cpu_we_i
  PIN gpio_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 296.000 267.630 300.000 ;
    END
  END gpio_ack_i
  PIN gpio_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 296.000 282.810 300.000 ;
    END
  END gpio_adr_o[0]
  PIN gpio_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 296.000 368.370 300.000 ;
    END
  END gpio_adr_o[10]
  PIN gpio_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 296.000 375.730 300.000 ;
    END
  END gpio_adr_o[11]
  PIN gpio_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 296.000 383.550 300.000 ;
    END
  END gpio_adr_o[12]
  PIN gpio_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 296.000 390.910 300.000 ;
    END
  END gpio_adr_o[13]
  PIN gpio_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 296.000 398.730 300.000 ;
    END
  END gpio_adr_o[14]
  PIN gpio_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 296.000 406.090 300.000 ;
    END
  END gpio_adr_o[15]
  PIN gpio_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 296.000 413.450 300.000 ;
    END
  END gpio_adr_o[16]
  PIN gpio_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 296.000 421.270 300.000 ;
    END
  END gpio_adr_o[17]
  PIN gpio_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 296.000 428.630 300.000 ;
    END
  END gpio_adr_o[18]
  PIN gpio_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 296.000 436.450 300.000 ;
    END
  END gpio_adr_o[19]
  PIN gpio_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 296.000 292.930 300.000 ;
    END
  END gpio_adr_o[1]
  PIN gpio_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 296.000 443.810 300.000 ;
    END
  END gpio_adr_o[20]
  PIN gpio_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 296.000 451.170 300.000 ;
    END
  END gpio_adr_o[21]
  PIN gpio_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.710 296.000 458.990 300.000 ;
    END
  END gpio_adr_o[22]
  PIN gpio_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 296.000 466.350 300.000 ;
    END
  END gpio_adr_o[23]
  PIN gpio_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 296.000 474.170 300.000 ;
    END
  END gpio_adr_o[24]
  PIN gpio_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.250 296.000 481.530 300.000 ;
    END
  END gpio_adr_o[25]
  PIN gpio_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 296.000 488.890 300.000 ;
    END
  END gpio_adr_o[26]
  PIN gpio_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 296.000 496.710 300.000 ;
    END
  END gpio_adr_o[27]
  PIN gpio_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 296.000 504.070 300.000 ;
    END
  END gpio_adr_o[28]
  PIN gpio_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 296.000 511.890 300.000 ;
    END
  END gpio_adr_o[29]
  PIN gpio_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 296.000 303.050 300.000 ;
    END
  END gpio_adr_o[2]
  PIN gpio_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 296.000 519.250 300.000 ;
    END
  END gpio_adr_o[30]
  PIN gpio_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 296.000 526.610 300.000 ;
    END
  END gpio_adr_o[31]
  PIN gpio_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 296.000 313.170 300.000 ;
    END
  END gpio_adr_o[3]
  PIN gpio_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 296.000 322.830 300.000 ;
    END
  END gpio_adr_o[4]
  PIN gpio_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 296.000 330.650 300.000 ;
    END
  END gpio_adr_o[5]
  PIN gpio_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 296.000 338.010 300.000 ;
    END
  END gpio_adr_o[6]
  PIN gpio_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 296.000 345.830 300.000 ;
    END
  END gpio_adr_o[7]
  PIN gpio_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 296.000 353.190 300.000 ;
    END
  END gpio_adr_o[8]
  PIN gpio_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 296.000 361.010 300.000 ;
    END
  END gpio_adr_o[9]
  PIN gpio_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 296.000 270.390 300.000 ;
    END
  END gpio_cyc_o
  PIN gpio_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 296.000 285.110 300.000 ;
    END
  END gpio_dat_i[0]
  PIN gpio_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 296.000 370.670 300.000 ;
    END
  END gpio_dat_i[10]
  PIN gpio_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 296.000 378.490 300.000 ;
    END
  END gpio_dat_i[11]
  PIN gpio_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 296.000 385.850 300.000 ;
    END
  END gpio_dat_i[12]
  PIN gpio_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 296.000 393.670 300.000 ;
    END
  END gpio_dat_i[13]
  PIN gpio_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 296.000 401.030 300.000 ;
    END
  END gpio_dat_i[14]
  PIN gpio_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 296.000 408.390 300.000 ;
    END
  END gpio_dat_i[15]
  PIN gpio_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 296.000 416.210 300.000 ;
    END
  END gpio_dat_i[16]
  PIN gpio_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 296.000 423.570 300.000 ;
    END
  END gpio_dat_i[17]
  PIN gpio_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.110 296.000 431.390 300.000 ;
    END
  END gpio_dat_i[18]
  PIN gpio_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 296.000 438.750 300.000 ;
    END
  END gpio_dat_i[19]
  PIN gpio_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 296.000 295.230 300.000 ;
    END
  END gpio_dat_i[1]
  PIN gpio_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 296.000 446.110 300.000 ;
    END
  END gpio_dat_i[20]
  PIN gpio_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 296.000 453.930 300.000 ;
    END
  END gpio_dat_i[21]
  PIN gpio_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 296.000 461.290 300.000 ;
    END
  END gpio_dat_i[22]
  PIN gpio_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.830 296.000 469.110 300.000 ;
    END
  END gpio_dat_i[23]
  PIN gpio_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 296.000 476.470 300.000 ;
    END
  END gpio_dat_i[24]
  PIN gpio_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 296.000 483.830 300.000 ;
    END
  END gpio_dat_i[25]
  PIN gpio_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 296.000 491.650 300.000 ;
    END
  END gpio_dat_i[26]
  PIN gpio_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 296.000 499.010 300.000 ;
    END
  END gpio_dat_i[27]
  PIN gpio_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 296.000 506.830 300.000 ;
    END
  END gpio_dat_i[28]
  PIN gpio_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 296.000 514.190 300.000 ;
    END
  END gpio_dat_i[29]
  PIN gpio_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 296.000 305.350 300.000 ;
    END
  END gpio_dat_i[2]
  PIN gpio_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 296.000 521.550 300.000 ;
    END
  END gpio_dat_i[30]
  PIN gpio_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 296.000 529.370 300.000 ;
    END
  END gpio_dat_i[31]
  PIN gpio_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 296.000 315.470 300.000 ;
    END
  END gpio_dat_i[3]
  PIN gpio_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 296.000 325.590 300.000 ;
    END
  END gpio_dat_i[4]
  PIN gpio_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 296.000 332.950 300.000 ;
    END
  END gpio_dat_i[5]
  PIN gpio_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 296.000 340.770 300.000 ;
    END
  END gpio_dat_i[6]
  PIN gpio_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 296.000 348.130 300.000 ;
    END
  END gpio_dat_i[7]
  PIN gpio_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 296.000 355.950 300.000 ;
    END
  END gpio_dat_i[8]
  PIN gpio_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 296.000 363.310 300.000 ;
    END
  END gpio_dat_i[9]
  PIN gpio_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 296.000 287.870 300.000 ;
    END
  END gpio_dat_o[0]
  PIN gpio_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 296.000 373.430 300.000 ;
    END
  END gpio_dat_o[10]
  PIN gpio_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 296.000 380.790 300.000 ;
    END
  END gpio_dat_o[11]
  PIN gpio_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 296.000 388.610 300.000 ;
    END
  END gpio_dat_o[12]
  PIN gpio_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 296.000 395.970 300.000 ;
    END
  END gpio_dat_o[13]
  PIN gpio_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 296.000 403.330 300.000 ;
    END
  END gpio_dat_o[14]
  PIN gpio_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 296.000 411.150 300.000 ;
    END
  END gpio_dat_o[15]
  PIN gpio_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 296.000 418.510 300.000 ;
    END
  END gpio_dat_o[16]
  PIN gpio_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 296.000 426.330 300.000 ;
    END
  END gpio_dat_o[17]
  PIN gpio_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 296.000 433.690 300.000 ;
    END
  END gpio_dat_o[18]
  PIN gpio_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 296.000 441.050 300.000 ;
    END
  END gpio_dat_o[19]
  PIN gpio_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 296.000 297.990 300.000 ;
    END
  END gpio_dat_o[1]
  PIN gpio_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 296.000 448.870 300.000 ;
    END
  END gpio_dat_o[20]
  PIN gpio_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 296.000 456.230 300.000 ;
    END
  END gpio_dat_o[21]
  PIN gpio_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 296.000 464.050 300.000 ;
    END
  END gpio_dat_o[22]
  PIN gpio_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 296.000 471.410 300.000 ;
    END
  END gpio_dat_o[23]
  PIN gpio_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 296.000 479.230 300.000 ;
    END
  END gpio_dat_o[24]
  PIN gpio_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 296.000 486.590 300.000 ;
    END
  END gpio_dat_o[25]
  PIN gpio_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.670 296.000 493.950 300.000 ;
    END
  END gpio_dat_o[26]
  PIN gpio_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.490 296.000 501.770 300.000 ;
    END
  END gpio_dat_o[27]
  PIN gpio_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 296.000 509.130 300.000 ;
    END
  END gpio_dat_o[28]
  PIN gpio_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 296.000 516.950 300.000 ;
    END
  END gpio_dat_o[29]
  PIN gpio_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 296.000 308.110 300.000 ;
    END
  END gpio_dat_o[2]
  PIN gpio_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 296.000 524.310 300.000 ;
    END
  END gpio_dat_o[30]
  PIN gpio_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 296.000 531.670 300.000 ;
    END
  END gpio_dat_o[31]
  PIN gpio_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 296.000 318.230 300.000 ;
    END
  END gpio_dat_o[3]
  PIN gpio_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 296.000 327.890 300.000 ;
    END
  END gpio_dat_o[4]
  PIN gpio_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 296.000 335.710 300.000 ;
    END
  END gpio_dat_o[5]
  PIN gpio_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 296.000 343.070 300.000 ;
    END
  END gpio_dat_o[6]
  PIN gpio_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 296.000 350.890 300.000 ;
    END
  END gpio_dat_o[7]
  PIN gpio_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 296.000 358.250 300.000 ;
    END
  END gpio_dat_o[8]
  PIN gpio_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 296.000 365.610 300.000 ;
    END
  END gpio_dat_o[9]
  PIN gpio_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 296.000 272.690 300.000 ;
    END
  END gpio_err_i
  PIN gpio_rty_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 296.000 275.450 300.000 ;
    END
  END gpio_rty_i
  PIN gpio_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 296.000 290.170 300.000 ;
    END
  END gpio_sel_o[0]
  PIN gpio_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 296.000 300.290 300.000 ;
    END
  END gpio_sel_o[1]
  PIN gpio_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 296.000 310.410 300.000 ;
    END
  END gpio_sel_o[2]
  PIN gpio_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 296.000 320.530 300.000 ;
    END
  END gpio_sel_o[3]
  PIN gpio_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 296.000 277.750 300.000 ;
    END
  END gpio_stb_o
  PIN gpio_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 296.000 280.510 300.000 ;
    END
  END gpio_we_o
  PIN ksc_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 296.000 534.430 300.000 ;
    END
  END ksc_ack_i
  PIN ksc_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 296.000 549.610 300.000 ;
    END
  END ksc_adr_o[0]
  PIN ksc_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 296.000 635.170 300.000 ;
    END
  END ksc_adr_o[10]
  PIN ksc_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.250 296.000 642.530 300.000 ;
    END
  END ksc_adr_o[11]
  PIN ksc_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 296.000 649.890 300.000 ;
    END
  END ksc_adr_o[12]
  PIN ksc_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 296.000 657.710 300.000 ;
    END
  END ksc_adr_o[13]
  PIN ksc_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.790 296.000 665.070 300.000 ;
    END
  END ksc_adr_o[14]
  PIN ksc_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 296.000 672.890 300.000 ;
    END
  END ksc_adr_o[15]
  PIN ksc_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 296.000 680.250 300.000 ;
    END
  END ksc_adr_o[16]
  PIN ksc_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 296.000 687.610 300.000 ;
    END
  END ksc_adr_o[17]
  PIN ksc_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.150 296.000 695.430 300.000 ;
    END
  END ksc_adr_o[18]
  PIN ksc_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 296.000 702.790 300.000 ;
    END
  END ksc_adr_o[19]
  PIN ksc_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 296.000 559.730 300.000 ;
    END
  END ksc_adr_o[1]
  PIN ksc_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 296.000 710.610 300.000 ;
    END
  END ksc_adr_o[20]
  PIN ksc_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 296.000 717.970 300.000 ;
    END
  END ksc_adr_o[21]
  PIN ksc_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 296.000 725.330 300.000 ;
    END
  END ksc_adr_o[22]
  PIN ksc_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 296.000 733.150 300.000 ;
    END
  END ksc_adr_o[23]
  PIN ksc_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.230 296.000 740.510 300.000 ;
    END
  END ksc_adr_o[24]
  PIN ksc_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 296.000 748.330 300.000 ;
    END
  END ksc_adr_o[25]
  PIN ksc_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.410 296.000 755.690 300.000 ;
    END
  END ksc_adr_o[26]
  PIN ksc_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.770 296.000 763.050 300.000 ;
    END
  END ksc_adr_o[27]
  PIN ksc_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.590 296.000 770.870 300.000 ;
    END
  END ksc_adr_o[28]
  PIN ksc_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 296.000 778.230 300.000 ;
    END
  END ksc_adr_o[29]
  PIN ksc_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.110 296.000 569.390 300.000 ;
    END
  END ksc_adr_o[2]
  PIN ksc_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 296.000 786.050 300.000 ;
    END
  END ksc_adr_o[30]
  PIN ksc_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 296.000 793.410 300.000 ;
    END
  END ksc_adr_o[31]
  PIN ksc_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 296.000 579.510 300.000 ;
    END
  END ksc_adr_o[3]
  PIN ksc_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 296.000 589.630 300.000 ;
    END
  END ksc_adr_o[4]
  PIN ksc_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.170 296.000 597.450 300.000 ;
    END
  END ksc_adr_o[5]
  PIN ksc_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 296.000 604.810 300.000 ;
    END
  END ksc_adr_o[6]
  PIN ksc_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 296.000 612.170 300.000 ;
    END
  END ksc_adr_o[7]
  PIN ksc_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 296.000 619.990 300.000 ;
    END
  END ksc_adr_o[8]
  PIN ksc_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.070 296.000 627.350 300.000 ;
    END
  END ksc_adr_o[9]
  PIN ksc_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 296.000 536.730 300.000 ;
    END
  END ksc_cyc_o
  PIN ksc_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 296.000 551.910 300.000 ;
    END
  END ksc_dat_i[0]
  PIN ksc_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 296.000 637.470 300.000 ;
    END
  END ksc_dat_i[10]
  PIN ksc_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.550 296.000 644.830 300.000 ;
    END
  END ksc_dat_i[11]
  PIN ksc_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 296.000 652.650 300.000 ;
    END
  END ksc_dat_i[12]
  PIN ksc_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.730 296.000 660.010 300.000 ;
    END
  END ksc_dat_i[13]
  PIN ksc_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 296.000 667.830 300.000 ;
    END
  END ksc_dat_i[14]
  PIN ksc_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 296.000 675.190 300.000 ;
    END
  END ksc_dat_i[15]
  PIN ksc_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.270 296.000 682.550 300.000 ;
    END
  END ksc_dat_i[16]
  PIN ksc_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 296.000 690.370 300.000 ;
    END
  END ksc_dat_i[17]
  PIN ksc_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 296.000 697.730 300.000 ;
    END
  END ksc_dat_i[18]
  PIN ksc_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 296.000 705.550 300.000 ;
    END
  END ksc_dat_i[19]
  PIN ksc_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 296.000 562.030 300.000 ;
    END
  END ksc_dat_i[1]
  PIN ksc_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 296.000 712.910 300.000 ;
    END
  END ksc_dat_i[20]
  PIN ksc_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 296.000 720.730 300.000 ;
    END
  END ksc_dat_i[21]
  PIN ksc_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 296.000 728.090 300.000 ;
    END
  END ksc_dat_i[22]
  PIN ksc_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 296.000 735.450 300.000 ;
    END
  END ksc_dat_i[23]
  PIN ksc_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.990 296.000 743.270 300.000 ;
    END
  END ksc_dat_i[24]
  PIN ksc_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 296.000 750.630 300.000 ;
    END
  END ksc_dat_i[25]
  PIN ksc_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 296.000 758.450 300.000 ;
    END
  END ksc_dat_i[26]
  PIN ksc_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 296.000 765.810 300.000 ;
    END
  END ksc_dat_i[27]
  PIN ksc_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 296.000 773.170 300.000 ;
    END
  END ksc_dat_i[28]
  PIN ksc_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.710 296.000 780.990 300.000 ;
    END
  END ksc_dat_i[29]
  PIN ksc_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.870 296.000 572.150 300.000 ;
    END
  END ksc_dat_i[2]
  PIN ksc_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.070 296.000 788.350 300.000 ;
    END
  END ksc_dat_i[30]
  PIN ksc_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 296.000 796.170 300.000 ;
    END
  END ksc_dat_i[31]
  PIN ksc_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 296.000 582.270 300.000 ;
    END
  END ksc_dat_i[3]
  PIN ksc_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 296.000 592.390 300.000 ;
    END
  END ksc_dat_i[4]
  PIN ksc_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 296.000 599.750 300.000 ;
    END
  END ksc_dat_i[5]
  PIN ksc_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.830 296.000 607.110 300.000 ;
    END
  END ksc_dat_i[6]
  PIN ksc_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 296.000 614.930 300.000 ;
    END
  END ksc_dat_i[7]
  PIN ksc_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.010 296.000 622.290 300.000 ;
    END
  END ksc_dat_i[8]
  PIN ksc_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 296.000 630.110 300.000 ;
    END
  END ksc_dat_i[9]
  PIN ksc_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 296.000 554.670 300.000 ;
    END
  END ksc_dat_o[0]
  PIN ksc_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.950 296.000 640.230 300.000 ;
    END
  END ksc_dat_o[10]
  PIN ksc_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 296.000 647.590 300.000 ;
    END
  END ksc_dat_o[11]
  PIN ksc_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.670 296.000 654.950 300.000 ;
    END
  END ksc_dat_o[12]
  PIN ksc_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 296.000 662.770 300.000 ;
    END
  END ksc_dat_o[13]
  PIN ksc_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 296.000 670.130 300.000 ;
    END
  END ksc_dat_o[14]
  PIN ksc_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.670 296.000 677.950 300.000 ;
    END
  END ksc_dat_o[15]
  PIN ksc_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 296.000 685.310 300.000 ;
    END
  END ksc_dat_o[16]
  PIN ksc_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 296.000 692.670 300.000 ;
    END
  END ksc_dat_o[17]
  PIN ksc_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 296.000 700.490 300.000 ;
    END
  END ksc_dat_o[18]
  PIN ksc_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 296.000 707.850 300.000 ;
    END
  END ksc_dat_o[19]
  PIN ksc_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 296.000 564.330 300.000 ;
    END
  END ksc_dat_o[1]
  PIN ksc_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 296.000 715.670 300.000 ;
    END
  END ksc_dat_o[20]
  PIN ksc_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.750 296.000 723.030 300.000 ;
    END
  END ksc_dat_o[21]
  PIN ksc_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 296.000 730.390 300.000 ;
    END
  END ksc_dat_o[22]
  PIN ksc_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 296.000 738.210 300.000 ;
    END
  END ksc_dat_o[23]
  PIN ksc_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 296.000 745.570 300.000 ;
    END
  END ksc_dat_o[24]
  PIN ksc_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.110 296.000 753.390 300.000 ;
    END
  END ksc_dat_o[25]
  PIN ksc_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.470 296.000 760.750 300.000 ;
    END
  END ksc_dat_o[26]
  PIN ksc_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 296.000 768.110 300.000 ;
    END
  END ksc_dat_o[27]
  PIN ksc_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 296.000 775.930 300.000 ;
    END
  END ksc_dat_o[28]
  PIN ksc_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 296.000 783.290 300.000 ;
    END
  END ksc_dat_o[29]
  PIN ksc_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 296.000 574.450 300.000 ;
    END
  END ksc_dat_o[2]
  PIN ksc_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.830 296.000 791.110 300.000 ;
    END
  END ksc_dat_o[30]
  PIN ksc_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 296.000 798.470 300.000 ;
    END
  END ksc_dat_o[31]
  PIN ksc_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 296.000 584.570 300.000 ;
    END
  END ksc_dat_o[3]
  PIN ksc_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 296.000 594.690 300.000 ;
    END
  END ksc_dat_o[4]
  PIN ksc_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.770 296.000 602.050 300.000 ;
    END
  END ksc_dat_o[5]
  PIN ksc_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 296.000 609.870 300.000 ;
    END
  END ksc_dat_o[6]
  PIN ksc_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.950 296.000 617.230 300.000 ;
    END
  END ksc_dat_o[7]
  PIN ksc_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 296.000 625.050 300.000 ;
    END
  END ksc_dat_o[8]
  PIN ksc_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 296.000 632.410 300.000 ;
    END
  END ksc_dat_o[9]
  PIN ksc_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 296.000 539.490 300.000 ;
    END
  END ksc_err_i
  PIN ksc_rty_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 296.000 541.790 300.000 ;
    END
  END ksc_rty_i
  PIN ksc_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 296.000 556.970 300.000 ;
    END
  END ksc_sel_o[0]
  PIN ksc_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 296.000 567.090 300.000 ;
    END
  END ksc_sel_o[1]
  PIN ksc_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 296.000 577.210 300.000 ;
    END
  END ksc_sel_o[2]
  PIN ksc_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 296.000 587.330 300.000 ;
    END
  END ksc_sel_o[3]
  PIN ksc_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 296.000 544.550 300.000 ;
    END
  END ksc_stb_o
  PIN ksc_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.570 296.000 546.850 300.000 ;
    END
  END ksc_we_o
  PIN spi_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 296.000 1.290 300.000 ;
    END
  END spi_ack_i
  PIN spi_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 296.000 16.010 300.000 ;
    END
  END spi_adr_o[0]
  PIN spi_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 296.000 101.570 300.000 ;
    END
  END spi_adr_o[10]
  PIN spi_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 296.000 109.390 300.000 ;
    END
  END spi_adr_o[11]
  PIN spi_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 296.000 116.750 300.000 ;
    END
  END spi_adr_o[12]
  PIN spi_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 296.000 124.110 300.000 ;
    END
  END spi_adr_o[13]
  PIN spi_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 296.000 131.930 300.000 ;
    END
  END spi_adr_o[14]
  PIN spi_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 296.000 139.290 300.000 ;
    END
  END spi_adr_o[15]
  PIN spi_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 296.000 147.110 300.000 ;
    END
  END spi_adr_o[16]
  PIN spi_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 296.000 154.470 300.000 ;
    END
  END spi_adr_o[17]
  PIN spi_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 296.000 161.830 300.000 ;
    END
  END spi_adr_o[18]
  PIN spi_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 296.000 169.650 300.000 ;
    END
  END spi_adr_o[19]
  PIN spi_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 296.000 26.130 300.000 ;
    END
  END spi_adr_o[1]
  PIN spi_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 296.000 177.010 300.000 ;
    END
  END spi_adr_o[20]
  PIN spi_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 296.000 184.830 300.000 ;
    END
  END spi_adr_o[21]
  PIN spi_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 296.000 192.190 300.000 ;
    END
  END spi_adr_o[22]
  PIN spi_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 296.000 200.010 300.000 ;
    END
  END spi_adr_o[23]
  PIN spi_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 296.000 207.370 300.000 ;
    END
  END spi_adr_o[24]
  PIN spi_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 296.000 214.730 300.000 ;
    END
  END spi_adr_o[25]
  PIN spi_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 296.000 222.550 300.000 ;
    END
  END spi_adr_o[26]
  PIN spi_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 296.000 229.910 300.000 ;
    END
  END spi_adr_o[27]
  PIN spi_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 296.000 237.730 300.000 ;
    END
  END spi_adr_o[28]
  PIN spi_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 296.000 245.090 300.000 ;
    END
  END spi_adr_o[29]
  PIN spi_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 296.000 36.250 300.000 ;
    END
  END spi_adr_o[2]
  PIN spi_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 296.000 252.450 300.000 ;
    END
  END spi_adr_o[30]
  PIN spi_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 296.000 260.270 300.000 ;
    END
  END spi_adr_o[31]
  PIN spi_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 296.000 46.370 300.000 ;
    END
  END spi_adr_o[3]
  PIN spi_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 296.000 56.490 300.000 ;
    END
  END spi_adr_o[4]
  PIN spi_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 296.000 63.850 300.000 ;
    END
  END spi_adr_o[5]
  PIN spi_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 296.000 71.670 300.000 ;
    END
  END spi_adr_o[6]
  PIN spi_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 296.000 79.030 300.000 ;
    END
  END spi_adr_o[7]
  PIN spi_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 296.000 86.390 300.000 ;
    END
  END spi_adr_o[8]
  PIN spi_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 296.000 94.210 300.000 ;
    END
  END spi_adr_o[9]
  PIN spi_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 296.000 3.590 300.000 ;
    END
  END spi_cyc_o
  PIN spi_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 296.000 18.770 300.000 ;
    END
  END spi_dat_i[0]
  PIN spi_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 296.000 104.330 300.000 ;
    END
  END spi_dat_i[10]
  PIN spi_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 296.000 111.690 300.000 ;
    END
  END spi_dat_i[11]
  PIN spi_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 296.000 119.510 300.000 ;
    END
  END spi_dat_i[12]
  PIN spi_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 296.000 126.870 300.000 ;
    END
  END spi_dat_i[13]
  PIN spi_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 296.000 134.230 300.000 ;
    END
  END spi_dat_i[14]
  PIN spi_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 296.000 142.050 300.000 ;
    END
  END spi_dat_i[15]
  PIN spi_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 296.000 149.410 300.000 ;
    END
  END spi_dat_i[16]
  PIN spi_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 296.000 157.230 300.000 ;
    END
  END spi_dat_i[17]
  PIN spi_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 296.000 164.590 300.000 ;
    END
  END spi_dat_i[18]
  PIN spi_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 296.000 171.950 300.000 ;
    END
  END spi_dat_i[19]
  PIN spi_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 296.000 28.890 300.000 ;
    END
  END spi_dat_i[1]
  PIN spi_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 296.000 179.770 300.000 ;
    END
  END spi_dat_i[20]
  PIN spi_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 296.000 187.130 300.000 ;
    END
  END spi_dat_i[21]
  PIN spi_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 296.000 194.950 300.000 ;
    END
  END spi_dat_i[22]
  PIN spi_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 296.000 202.310 300.000 ;
    END
  END spi_dat_i[23]
  PIN spi_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 296.000 209.670 300.000 ;
    END
  END spi_dat_i[24]
  PIN spi_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 296.000 217.490 300.000 ;
    END
  END spi_dat_i[25]
  PIN spi_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 296.000 224.850 300.000 ;
    END
  END spi_dat_i[26]
  PIN spi_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 296.000 232.670 300.000 ;
    END
  END spi_dat_i[27]
  PIN spi_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 296.000 240.030 300.000 ;
    END
  END spi_dat_i[28]
  PIN spi_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 296.000 247.390 300.000 ;
    END
  END spi_dat_i[29]
  PIN spi_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 296.000 39.010 300.000 ;
    END
  END spi_dat_i[2]
  PIN spi_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 296.000 255.210 300.000 ;
    END
  END spi_dat_i[30]
  PIN spi_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 296.000 262.570 300.000 ;
    END
  END spi_dat_i[31]
  PIN spi_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 296.000 48.670 300.000 ;
    END
  END spi_dat_i[3]
  PIN spi_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 296.000 58.790 300.000 ;
    END
  END spi_dat_i[4]
  PIN spi_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 296.000 66.610 300.000 ;
    END
  END spi_dat_i[5]
  PIN spi_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 296.000 73.970 300.000 ;
    END
  END spi_dat_i[6]
  PIN spi_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 296.000 81.330 300.000 ;
    END
  END spi_dat_i[7]
  PIN spi_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 296.000 89.150 300.000 ;
    END
  END spi_dat_i[8]
  PIN spi_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 296.000 96.510 300.000 ;
    END
  END spi_dat_i[9]
  PIN spi_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 296.000 21.070 300.000 ;
    END
  END spi_dat_o[0]
  PIN spi_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 296.000 106.630 300.000 ;
    END
  END spi_dat_o[10]
  PIN spi_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 296.000 114.450 300.000 ;
    END
  END spi_dat_o[11]
  PIN spi_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 296.000 121.810 300.000 ;
    END
  END spi_dat_o[12]
  PIN spi_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 296.000 129.170 300.000 ;
    END
  END spi_dat_o[13]
  PIN spi_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 296.000 136.990 300.000 ;
    END
  END spi_dat_o[14]
  PIN spi_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 296.000 144.350 300.000 ;
    END
  END spi_dat_o[15]
  PIN spi_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 296.000 152.170 300.000 ;
    END
  END spi_dat_o[16]
  PIN spi_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 296.000 159.530 300.000 ;
    END
  END spi_dat_o[17]
  PIN spi_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 296.000 166.890 300.000 ;
    END
  END spi_dat_o[18]
  PIN spi_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 296.000 174.710 300.000 ;
    END
  END spi_dat_o[19]
  PIN spi_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 296.000 31.190 300.000 ;
    END
  END spi_dat_o[1]
  PIN spi_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 296.000 182.070 300.000 ;
    END
  END spi_dat_o[20]
  PIN spi_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 296.000 189.890 300.000 ;
    END
  END spi_dat_o[21]
  PIN spi_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 296.000 197.250 300.000 ;
    END
  END spi_dat_o[22]
  PIN spi_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 296.000 204.610 300.000 ;
    END
  END spi_dat_o[23]
  PIN spi_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 296.000 212.430 300.000 ;
    END
  END spi_dat_o[24]
  PIN spi_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 296.000 219.790 300.000 ;
    END
  END spi_dat_o[25]
  PIN spi_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 296.000 227.610 300.000 ;
    END
  END spi_dat_o[26]
  PIN spi_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 296.000 234.970 300.000 ;
    END
  END spi_dat_o[27]
  PIN spi_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 296.000 242.330 300.000 ;
    END
  END spi_dat_o[28]
  PIN spi_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 296.000 250.150 300.000 ;
    END
  END spi_dat_o[29]
  PIN spi_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 296.000 41.310 300.000 ;
    END
  END spi_dat_o[2]
  PIN spi_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 296.000 257.510 300.000 ;
    END
  END spi_dat_o[30]
  PIN spi_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 296.000 265.330 300.000 ;
    END
  END spi_dat_o[31]
  PIN spi_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 296.000 51.430 300.000 ;
    END
  END spi_dat_o[3]
  PIN spi_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 296.000 61.550 300.000 ;
    END
  END spi_dat_o[4]
  PIN spi_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 296.000 68.910 300.000 ;
    END
  END spi_dat_o[5]
  PIN spi_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 296.000 76.730 300.000 ;
    END
  END spi_dat_o[6]
  PIN spi_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 296.000 84.090 300.000 ;
    END
  END spi_dat_o[7]
  PIN spi_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 296.000 91.450 300.000 ;
    END
  END spi_dat_o[8]
  PIN spi_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 296.000 99.270 300.000 ;
    END
  END spi_dat_o[9]
  PIN spi_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 296.000 5.890 300.000 ;
    END
  END spi_err_i
  PIN spi_rty_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 296.000 8.650 300.000 ;
    END
  END spi_rty_i
  PIN spi_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 296.000 23.830 300.000 ;
    END
  END spi_sel_o[0]
  PIN spi_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 296.000 33.950 300.000 ;
    END
  END spi_sel_o[1]
  PIN spi_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 296.000 43.610 300.000 ;
    END
  END spi_sel_o[2]
  PIN spi_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 296.000 53.730 300.000 ;
    END
  END spi_sel_o[3]
  PIN spi_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 296.000 10.950 300.000 ;
    END
  END spi_stb_o
  PIN spi_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 296.000 13.710 300.000 ;
    END
  END spi_we_o
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 288.560 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 794.420 288.405 ;
      LAYER met1 ;
        RECT 0.990 6.500 796.190 296.100 ;
      LAYER met2 ;
        RECT 1.570 295.720 3.030 299.725 ;
        RECT 3.870 295.720 5.330 299.725 ;
        RECT 6.170 295.720 8.090 299.725 ;
        RECT 8.930 295.720 10.390 299.725 ;
        RECT 11.230 295.720 13.150 299.725 ;
        RECT 13.990 295.720 15.450 299.725 ;
        RECT 16.290 295.720 18.210 299.725 ;
        RECT 19.050 295.720 20.510 299.725 ;
        RECT 21.350 295.720 23.270 299.725 ;
        RECT 24.110 295.720 25.570 299.725 ;
        RECT 26.410 295.720 28.330 299.725 ;
        RECT 29.170 295.720 30.630 299.725 ;
        RECT 31.470 295.720 33.390 299.725 ;
        RECT 34.230 295.720 35.690 299.725 ;
        RECT 36.530 295.720 38.450 299.725 ;
        RECT 39.290 295.720 40.750 299.725 ;
        RECT 41.590 295.720 43.050 299.725 ;
        RECT 43.890 295.720 45.810 299.725 ;
        RECT 46.650 295.720 48.110 299.725 ;
        RECT 48.950 295.720 50.870 299.725 ;
        RECT 51.710 295.720 53.170 299.725 ;
        RECT 54.010 295.720 55.930 299.725 ;
        RECT 56.770 295.720 58.230 299.725 ;
        RECT 59.070 295.720 60.990 299.725 ;
        RECT 61.830 295.720 63.290 299.725 ;
        RECT 64.130 295.720 66.050 299.725 ;
        RECT 66.890 295.720 68.350 299.725 ;
        RECT 69.190 295.720 71.110 299.725 ;
        RECT 71.950 295.720 73.410 299.725 ;
        RECT 74.250 295.720 76.170 299.725 ;
        RECT 77.010 295.720 78.470 299.725 ;
        RECT 79.310 295.720 80.770 299.725 ;
        RECT 81.610 295.720 83.530 299.725 ;
        RECT 84.370 295.720 85.830 299.725 ;
        RECT 86.670 295.720 88.590 299.725 ;
        RECT 89.430 295.720 90.890 299.725 ;
        RECT 91.730 295.720 93.650 299.725 ;
        RECT 94.490 295.720 95.950 299.725 ;
        RECT 96.790 295.720 98.710 299.725 ;
        RECT 99.550 295.720 101.010 299.725 ;
        RECT 101.850 295.720 103.770 299.725 ;
        RECT 104.610 295.720 106.070 299.725 ;
        RECT 106.910 295.720 108.830 299.725 ;
        RECT 109.670 295.720 111.130 299.725 ;
        RECT 111.970 295.720 113.890 299.725 ;
        RECT 114.730 295.720 116.190 299.725 ;
        RECT 117.030 295.720 118.950 299.725 ;
        RECT 119.790 295.720 121.250 299.725 ;
        RECT 122.090 295.720 123.550 299.725 ;
        RECT 124.390 295.720 126.310 299.725 ;
        RECT 127.150 295.720 128.610 299.725 ;
        RECT 129.450 295.720 131.370 299.725 ;
        RECT 132.210 295.720 133.670 299.725 ;
        RECT 134.510 295.720 136.430 299.725 ;
        RECT 137.270 295.720 138.730 299.725 ;
        RECT 139.570 295.720 141.490 299.725 ;
        RECT 142.330 295.720 143.790 299.725 ;
        RECT 144.630 295.720 146.550 299.725 ;
        RECT 147.390 295.720 148.850 299.725 ;
        RECT 149.690 295.720 151.610 299.725 ;
        RECT 152.450 295.720 153.910 299.725 ;
        RECT 154.750 295.720 156.670 299.725 ;
        RECT 157.510 295.720 158.970 299.725 ;
        RECT 159.810 295.720 161.270 299.725 ;
        RECT 162.110 295.720 164.030 299.725 ;
        RECT 164.870 295.720 166.330 299.725 ;
        RECT 167.170 295.720 169.090 299.725 ;
        RECT 169.930 295.720 171.390 299.725 ;
        RECT 172.230 295.720 174.150 299.725 ;
        RECT 174.990 295.720 176.450 299.725 ;
        RECT 177.290 295.720 179.210 299.725 ;
        RECT 180.050 295.720 181.510 299.725 ;
        RECT 182.350 295.720 184.270 299.725 ;
        RECT 185.110 295.720 186.570 299.725 ;
        RECT 187.410 295.720 189.330 299.725 ;
        RECT 190.170 295.720 191.630 299.725 ;
        RECT 192.470 295.720 194.390 299.725 ;
        RECT 195.230 295.720 196.690 299.725 ;
        RECT 197.530 295.720 199.450 299.725 ;
        RECT 200.290 295.720 201.750 299.725 ;
        RECT 202.590 295.720 204.050 299.725 ;
        RECT 204.890 295.720 206.810 299.725 ;
        RECT 207.650 295.720 209.110 299.725 ;
        RECT 209.950 295.720 211.870 299.725 ;
        RECT 212.710 295.720 214.170 299.725 ;
        RECT 215.010 295.720 216.930 299.725 ;
        RECT 217.770 295.720 219.230 299.725 ;
        RECT 220.070 295.720 221.990 299.725 ;
        RECT 222.830 295.720 224.290 299.725 ;
        RECT 225.130 295.720 227.050 299.725 ;
        RECT 227.890 295.720 229.350 299.725 ;
        RECT 230.190 295.720 232.110 299.725 ;
        RECT 232.950 295.720 234.410 299.725 ;
        RECT 235.250 295.720 237.170 299.725 ;
        RECT 238.010 295.720 239.470 299.725 ;
        RECT 240.310 295.720 241.770 299.725 ;
        RECT 242.610 295.720 244.530 299.725 ;
        RECT 245.370 295.720 246.830 299.725 ;
        RECT 247.670 295.720 249.590 299.725 ;
        RECT 250.430 295.720 251.890 299.725 ;
        RECT 252.730 295.720 254.650 299.725 ;
        RECT 255.490 295.720 256.950 299.725 ;
        RECT 257.790 295.720 259.710 299.725 ;
        RECT 260.550 295.720 262.010 299.725 ;
        RECT 262.850 295.720 264.770 299.725 ;
        RECT 265.610 295.720 267.070 299.725 ;
        RECT 267.910 295.720 269.830 299.725 ;
        RECT 270.670 295.720 272.130 299.725 ;
        RECT 272.970 295.720 274.890 299.725 ;
        RECT 275.730 295.720 277.190 299.725 ;
        RECT 278.030 295.720 279.950 299.725 ;
        RECT 280.790 295.720 282.250 299.725 ;
        RECT 283.090 295.720 284.550 299.725 ;
        RECT 285.390 295.720 287.310 299.725 ;
        RECT 288.150 295.720 289.610 299.725 ;
        RECT 290.450 295.720 292.370 299.725 ;
        RECT 293.210 295.720 294.670 299.725 ;
        RECT 295.510 295.720 297.430 299.725 ;
        RECT 298.270 295.720 299.730 299.725 ;
        RECT 300.570 295.720 302.490 299.725 ;
        RECT 303.330 295.720 304.790 299.725 ;
        RECT 305.630 295.720 307.550 299.725 ;
        RECT 308.390 295.720 309.850 299.725 ;
        RECT 310.690 295.720 312.610 299.725 ;
        RECT 313.450 295.720 314.910 299.725 ;
        RECT 315.750 295.720 317.670 299.725 ;
        RECT 318.510 295.720 319.970 299.725 ;
        RECT 320.810 295.720 322.270 299.725 ;
        RECT 323.110 295.720 325.030 299.725 ;
        RECT 325.870 295.720 327.330 299.725 ;
        RECT 328.170 295.720 330.090 299.725 ;
        RECT 330.930 295.720 332.390 299.725 ;
        RECT 333.230 295.720 335.150 299.725 ;
        RECT 335.990 295.720 337.450 299.725 ;
        RECT 338.290 295.720 340.210 299.725 ;
        RECT 341.050 295.720 342.510 299.725 ;
        RECT 343.350 295.720 345.270 299.725 ;
        RECT 346.110 295.720 347.570 299.725 ;
        RECT 348.410 295.720 350.330 299.725 ;
        RECT 351.170 295.720 352.630 299.725 ;
        RECT 353.470 295.720 355.390 299.725 ;
        RECT 356.230 295.720 357.690 299.725 ;
        RECT 358.530 295.720 360.450 299.725 ;
        RECT 361.290 295.720 362.750 299.725 ;
        RECT 363.590 295.720 365.050 299.725 ;
        RECT 365.890 295.720 367.810 299.725 ;
        RECT 368.650 295.720 370.110 299.725 ;
        RECT 370.950 295.720 372.870 299.725 ;
        RECT 373.710 295.720 375.170 299.725 ;
        RECT 376.010 295.720 377.930 299.725 ;
        RECT 378.770 295.720 380.230 299.725 ;
        RECT 381.070 295.720 382.990 299.725 ;
        RECT 383.830 295.720 385.290 299.725 ;
        RECT 386.130 295.720 388.050 299.725 ;
        RECT 388.890 295.720 390.350 299.725 ;
        RECT 391.190 295.720 393.110 299.725 ;
        RECT 393.950 295.720 395.410 299.725 ;
        RECT 396.250 295.720 398.170 299.725 ;
        RECT 399.010 295.720 400.470 299.725 ;
        RECT 401.310 295.720 402.770 299.725 ;
        RECT 403.610 295.720 405.530 299.725 ;
        RECT 406.370 295.720 407.830 299.725 ;
        RECT 408.670 295.720 410.590 299.725 ;
        RECT 411.430 295.720 412.890 299.725 ;
        RECT 413.730 295.720 415.650 299.725 ;
        RECT 416.490 295.720 417.950 299.725 ;
        RECT 418.790 295.720 420.710 299.725 ;
        RECT 421.550 295.720 423.010 299.725 ;
        RECT 423.850 295.720 425.770 299.725 ;
        RECT 426.610 295.720 428.070 299.725 ;
        RECT 428.910 295.720 430.830 299.725 ;
        RECT 431.670 295.720 433.130 299.725 ;
        RECT 433.970 295.720 435.890 299.725 ;
        RECT 436.730 295.720 438.190 299.725 ;
        RECT 439.030 295.720 440.490 299.725 ;
        RECT 441.330 295.720 443.250 299.725 ;
        RECT 444.090 295.720 445.550 299.725 ;
        RECT 446.390 295.720 448.310 299.725 ;
        RECT 449.150 295.720 450.610 299.725 ;
        RECT 451.450 295.720 453.370 299.725 ;
        RECT 454.210 295.720 455.670 299.725 ;
        RECT 456.510 295.720 458.430 299.725 ;
        RECT 459.270 295.720 460.730 299.725 ;
        RECT 461.570 295.720 463.490 299.725 ;
        RECT 464.330 295.720 465.790 299.725 ;
        RECT 466.630 295.720 468.550 299.725 ;
        RECT 469.390 295.720 470.850 299.725 ;
        RECT 471.690 295.720 473.610 299.725 ;
        RECT 474.450 295.720 475.910 299.725 ;
        RECT 476.750 295.720 478.670 299.725 ;
        RECT 479.510 295.720 480.970 299.725 ;
        RECT 481.810 295.720 483.270 299.725 ;
        RECT 484.110 295.720 486.030 299.725 ;
        RECT 486.870 295.720 488.330 299.725 ;
        RECT 489.170 295.720 491.090 299.725 ;
        RECT 491.930 295.720 493.390 299.725 ;
        RECT 494.230 295.720 496.150 299.725 ;
        RECT 496.990 295.720 498.450 299.725 ;
        RECT 499.290 295.720 501.210 299.725 ;
        RECT 502.050 295.720 503.510 299.725 ;
        RECT 504.350 295.720 506.270 299.725 ;
        RECT 507.110 295.720 508.570 299.725 ;
        RECT 509.410 295.720 511.330 299.725 ;
        RECT 512.170 295.720 513.630 299.725 ;
        RECT 514.470 295.720 516.390 299.725 ;
        RECT 517.230 295.720 518.690 299.725 ;
        RECT 519.530 295.720 520.990 299.725 ;
        RECT 521.830 295.720 523.750 299.725 ;
        RECT 524.590 295.720 526.050 299.725 ;
        RECT 526.890 295.720 528.810 299.725 ;
        RECT 529.650 295.720 531.110 299.725 ;
        RECT 531.950 295.720 533.870 299.725 ;
        RECT 534.710 295.720 536.170 299.725 ;
        RECT 537.010 295.720 538.930 299.725 ;
        RECT 539.770 295.720 541.230 299.725 ;
        RECT 542.070 295.720 543.990 299.725 ;
        RECT 544.830 295.720 546.290 299.725 ;
        RECT 547.130 295.720 549.050 299.725 ;
        RECT 549.890 295.720 551.350 299.725 ;
        RECT 552.190 295.720 554.110 299.725 ;
        RECT 554.950 295.720 556.410 299.725 ;
        RECT 557.250 295.720 559.170 299.725 ;
        RECT 560.010 295.720 561.470 299.725 ;
        RECT 562.310 295.720 563.770 299.725 ;
        RECT 564.610 295.720 566.530 299.725 ;
        RECT 567.370 295.720 568.830 299.725 ;
        RECT 569.670 295.720 571.590 299.725 ;
        RECT 572.430 295.720 573.890 299.725 ;
        RECT 574.730 295.720 576.650 299.725 ;
        RECT 577.490 295.720 578.950 299.725 ;
        RECT 579.790 295.720 581.710 299.725 ;
        RECT 582.550 295.720 584.010 299.725 ;
        RECT 584.850 295.720 586.770 299.725 ;
        RECT 587.610 295.720 589.070 299.725 ;
        RECT 589.910 295.720 591.830 299.725 ;
        RECT 592.670 295.720 594.130 299.725 ;
        RECT 594.970 295.720 596.890 299.725 ;
        RECT 597.730 295.720 599.190 299.725 ;
        RECT 600.030 295.720 601.490 299.725 ;
        RECT 602.330 295.720 604.250 299.725 ;
        RECT 605.090 295.720 606.550 299.725 ;
        RECT 607.390 295.720 609.310 299.725 ;
        RECT 610.150 295.720 611.610 299.725 ;
        RECT 612.450 295.720 614.370 299.725 ;
        RECT 615.210 295.720 616.670 299.725 ;
        RECT 617.510 295.720 619.430 299.725 ;
        RECT 620.270 295.720 621.730 299.725 ;
        RECT 622.570 295.720 624.490 299.725 ;
        RECT 625.330 295.720 626.790 299.725 ;
        RECT 627.630 295.720 629.550 299.725 ;
        RECT 630.390 295.720 631.850 299.725 ;
        RECT 632.690 295.720 634.610 299.725 ;
        RECT 635.450 295.720 636.910 299.725 ;
        RECT 637.750 295.720 639.670 299.725 ;
        RECT 640.510 295.720 641.970 299.725 ;
        RECT 642.810 295.720 644.270 299.725 ;
        RECT 645.110 295.720 647.030 299.725 ;
        RECT 647.870 295.720 649.330 299.725 ;
        RECT 650.170 295.720 652.090 299.725 ;
        RECT 652.930 295.720 654.390 299.725 ;
        RECT 655.230 295.720 657.150 299.725 ;
        RECT 657.990 295.720 659.450 299.725 ;
        RECT 660.290 295.720 662.210 299.725 ;
        RECT 663.050 295.720 664.510 299.725 ;
        RECT 665.350 295.720 667.270 299.725 ;
        RECT 668.110 295.720 669.570 299.725 ;
        RECT 670.410 295.720 672.330 299.725 ;
        RECT 673.170 295.720 674.630 299.725 ;
        RECT 675.470 295.720 677.390 299.725 ;
        RECT 678.230 295.720 679.690 299.725 ;
        RECT 680.530 295.720 681.990 299.725 ;
        RECT 682.830 295.720 684.750 299.725 ;
        RECT 685.590 295.720 687.050 299.725 ;
        RECT 687.890 295.720 689.810 299.725 ;
        RECT 690.650 295.720 692.110 299.725 ;
        RECT 692.950 295.720 694.870 299.725 ;
        RECT 695.710 295.720 697.170 299.725 ;
        RECT 698.010 295.720 699.930 299.725 ;
        RECT 700.770 295.720 702.230 299.725 ;
        RECT 703.070 295.720 704.990 299.725 ;
        RECT 705.830 295.720 707.290 299.725 ;
        RECT 708.130 295.720 710.050 299.725 ;
        RECT 710.890 295.720 712.350 299.725 ;
        RECT 713.190 295.720 715.110 299.725 ;
        RECT 715.950 295.720 717.410 299.725 ;
        RECT 718.250 295.720 720.170 299.725 ;
        RECT 721.010 295.720 722.470 299.725 ;
        RECT 723.310 295.720 724.770 299.725 ;
        RECT 725.610 295.720 727.530 299.725 ;
        RECT 728.370 295.720 729.830 299.725 ;
        RECT 730.670 295.720 732.590 299.725 ;
        RECT 733.430 295.720 734.890 299.725 ;
        RECT 735.730 295.720 737.650 299.725 ;
        RECT 738.490 295.720 739.950 299.725 ;
        RECT 740.790 295.720 742.710 299.725 ;
        RECT 743.550 295.720 745.010 299.725 ;
        RECT 745.850 295.720 747.770 299.725 ;
        RECT 748.610 295.720 750.070 299.725 ;
        RECT 750.910 295.720 752.830 299.725 ;
        RECT 753.670 295.720 755.130 299.725 ;
        RECT 755.970 295.720 757.890 299.725 ;
        RECT 758.730 295.720 760.190 299.725 ;
        RECT 761.030 295.720 762.490 299.725 ;
        RECT 763.330 295.720 765.250 299.725 ;
        RECT 766.090 295.720 767.550 299.725 ;
        RECT 768.390 295.720 770.310 299.725 ;
        RECT 771.150 295.720 772.610 299.725 ;
        RECT 773.450 295.720 775.370 299.725 ;
        RECT 776.210 295.720 777.670 299.725 ;
        RECT 778.510 295.720 780.430 299.725 ;
        RECT 781.270 295.720 782.730 299.725 ;
        RECT 783.570 295.720 785.490 299.725 ;
        RECT 786.330 295.720 787.790 299.725 ;
        RECT 788.630 295.720 790.550 299.725 ;
        RECT 791.390 295.720 792.850 299.725 ;
        RECT 793.690 295.720 795.610 299.725 ;
        RECT 796.450 295.720 797.910 299.725 ;
        RECT 1.020 1.515 798.400 295.720 ;
      LAYER met3 ;
        RECT 4.000 298.880 790.640 299.705 ;
        RECT 4.400 297.480 790.640 298.880 ;
        RECT 4.000 296.160 790.640 297.480 ;
        RECT 4.400 294.760 790.640 296.160 ;
        RECT 4.000 293.440 790.640 294.760 ;
        RECT 4.400 292.040 790.640 293.440 ;
        RECT 4.000 290.720 790.640 292.040 ;
        RECT 4.400 289.320 790.640 290.720 ;
        RECT 4.000 288.000 790.640 289.320 ;
        RECT 4.400 286.600 790.640 288.000 ;
        RECT 4.000 285.280 790.640 286.600 ;
        RECT 4.400 283.880 790.640 285.280 ;
        RECT 4.000 282.560 790.640 283.880 ;
        RECT 4.400 281.160 790.640 282.560 ;
        RECT 4.000 279.840 790.640 281.160 ;
        RECT 4.400 278.440 790.640 279.840 ;
        RECT 4.000 277.120 790.640 278.440 ;
        RECT 4.400 275.720 790.640 277.120 ;
        RECT 4.000 274.400 790.640 275.720 ;
        RECT 4.400 273.000 790.640 274.400 ;
        RECT 4.000 271.680 790.640 273.000 ;
        RECT 4.400 270.280 790.640 271.680 ;
        RECT 4.000 268.960 790.640 270.280 ;
        RECT 4.400 267.560 790.640 268.960 ;
        RECT 4.000 265.560 790.640 267.560 ;
        RECT 4.400 264.160 790.640 265.560 ;
        RECT 4.000 262.840 790.640 264.160 ;
        RECT 4.400 261.440 790.640 262.840 ;
        RECT 4.000 260.120 790.640 261.440 ;
        RECT 4.400 258.720 790.640 260.120 ;
        RECT 4.000 257.400 790.640 258.720 ;
        RECT 4.400 256.000 790.640 257.400 ;
        RECT 4.000 254.680 790.640 256.000 ;
        RECT 4.400 253.280 790.640 254.680 ;
        RECT 4.000 251.960 790.640 253.280 ;
        RECT 4.400 250.560 790.640 251.960 ;
        RECT 4.000 249.240 790.640 250.560 ;
        RECT 4.400 247.840 790.640 249.240 ;
        RECT 4.000 246.520 790.640 247.840 ;
        RECT 4.400 245.120 790.640 246.520 ;
        RECT 4.000 243.800 790.640 245.120 ;
        RECT 4.400 242.400 790.640 243.800 ;
        RECT 4.000 241.080 790.640 242.400 ;
        RECT 4.400 239.680 790.640 241.080 ;
        RECT 4.000 238.360 790.640 239.680 ;
        RECT 4.400 236.960 790.640 238.360 ;
        RECT 4.000 235.640 790.640 236.960 ;
        RECT 4.400 234.240 790.640 235.640 ;
        RECT 4.000 232.240 790.640 234.240 ;
        RECT 4.400 230.840 790.640 232.240 ;
        RECT 4.000 229.520 790.640 230.840 ;
        RECT 4.400 228.120 790.640 229.520 ;
        RECT 4.000 226.800 790.640 228.120 ;
        RECT 4.400 225.400 790.640 226.800 ;
        RECT 4.000 224.080 790.640 225.400 ;
        RECT 4.400 222.680 790.640 224.080 ;
        RECT 4.000 221.360 790.640 222.680 ;
        RECT 4.400 219.960 790.640 221.360 ;
        RECT 4.000 218.640 790.640 219.960 ;
        RECT 4.400 217.240 790.640 218.640 ;
        RECT 4.000 215.920 790.640 217.240 ;
        RECT 4.400 214.520 790.640 215.920 ;
        RECT 4.000 213.200 790.640 214.520 ;
        RECT 4.400 211.800 790.640 213.200 ;
        RECT 4.000 210.480 790.640 211.800 ;
        RECT 4.400 209.080 790.640 210.480 ;
        RECT 4.000 207.760 790.640 209.080 ;
        RECT 4.400 206.360 790.640 207.760 ;
        RECT 4.000 205.040 790.640 206.360 ;
        RECT 4.400 203.640 790.640 205.040 ;
        RECT 4.000 202.320 790.640 203.640 ;
        RECT 4.400 200.920 790.640 202.320 ;
        RECT 4.000 198.920 790.640 200.920 ;
        RECT 4.400 197.520 790.640 198.920 ;
        RECT 4.000 196.200 790.640 197.520 ;
        RECT 4.400 194.800 790.640 196.200 ;
        RECT 4.000 193.480 790.640 194.800 ;
        RECT 4.400 192.080 790.640 193.480 ;
        RECT 4.000 190.760 790.640 192.080 ;
        RECT 4.400 189.360 790.640 190.760 ;
        RECT 4.000 188.040 790.640 189.360 ;
        RECT 4.400 186.640 790.640 188.040 ;
        RECT 4.000 185.320 790.640 186.640 ;
        RECT 4.400 183.920 790.640 185.320 ;
        RECT 4.000 182.600 790.640 183.920 ;
        RECT 4.400 181.200 790.640 182.600 ;
        RECT 4.000 179.880 790.640 181.200 ;
        RECT 4.400 178.480 790.640 179.880 ;
        RECT 4.000 177.160 790.640 178.480 ;
        RECT 4.400 175.760 790.640 177.160 ;
        RECT 4.000 174.440 790.640 175.760 ;
        RECT 4.400 173.040 790.640 174.440 ;
        RECT 4.000 171.720 790.640 173.040 ;
        RECT 4.400 170.320 790.640 171.720 ;
        RECT 4.000 169.000 790.640 170.320 ;
        RECT 4.400 167.600 790.640 169.000 ;
        RECT 4.000 165.600 790.640 167.600 ;
        RECT 4.400 164.200 790.640 165.600 ;
        RECT 4.000 162.880 790.640 164.200 ;
        RECT 4.400 161.480 790.640 162.880 ;
        RECT 4.000 160.160 790.640 161.480 ;
        RECT 4.400 158.760 790.640 160.160 ;
        RECT 4.000 157.440 790.640 158.760 ;
        RECT 4.400 156.040 790.640 157.440 ;
        RECT 4.000 154.720 790.640 156.040 ;
        RECT 4.400 153.320 790.640 154.720 ;
        RECT 4.000 152.000 790.640 153.320 ;
        RECT 4.400 150.600 790.640 152.000 ;
        RECT 4.000 149.280 790.640 150.600 ;
        RECT 4.400 147.880 790.640 149.280 ;
        RECT 4.000 146.560 790.640 147.880 ;
        RECT 4.400 145.160 790.640 146.560 ;
        RECT 4.000 143.840 790.640 145.160 ;
        RECT 4.400 142.440 790.640 143.840 ;
        RECT 4.000 141.120 790.640 142.440 ;
        RECT 4.400 139.720 790.640 141.120 ;
        RECT 4.000 138.400 790.640 139.720 ;
        RECT 4.400 137.000 790.640 138.400 ;
        RECT 4.000 135.680 790.640 137.000 ;
        RECT 4.400 134.280 790.640 135.680 ;
        RECT 4.000 132.280 790.640 134.280 ;
        RECT 4.400 130.880 790.640 132.280 ;
        RECT 4.000 129.560 790.640 130.880 ;
        RECT 4.400 128.160 790.640 129.560 ;
        RECT 4.000 126.840 790.640 128.160 ;
        RECT 4.400 125.440 790.640 126.840 ;
        RECT 4.000 124.120 790.640 125.440 ;
        RECT 4.400 122.720 790.640 124.120 ;
        RECT 4.000 121.400 790.640 122.720 ;
        RECT 4.400 120.000 790.640 121.400 ;
        RECT 4.000 118.680 790.640 120.000 ;
        RECT 4.400 117.280 790.640 118.680 ;
        RECT 4.000 115.960 790.640 117.280 ;
        RECT 4.400 114.560 790.640 115.960 ;
        RECT 4.000 113.240 790.640 114.560 ;
        RECT 4.400 111.840 790.640 113.240 ;
        RECT 4.000 110.520 790.640 111.840 ;
        RECT 4.400 109.120 790.640 110.520 ;
        RECT 4.000 107.800 790.640 109.120 ;
        RECT 4.400 106.400 790.640 107.800 ;
        RECT 4.000 105.080 790.640 106.400 ;
        RECT 4.400 103.680 790.640 105.080 ;
        RECT 4.000 102.360 790.640 103.680 ;
        RECT 4.400 100.960 790.640 102.360 ;
        RECT 4.000 98.960 790.640 100.960 ;
        RECT 4.400 97.560 790.640 98.960 ;
        RECT 4.000 96.240 790.640 97.560 ;
        RECT 4.400 94.840 790.640 96.240 ;
        RECT 4.000 93.520 790.640 94.840 ;
        RECT 4.400 92.120 790.640 93.520 ;
        RECT 4.000 90.800 790.640 92.120 ;
        RECT 4.400 89.400 790.640 90.800 ;
        RECT 4.000 88.080 790.640 89.400 ;
        RECT 4.400 86.680 790.640 88.080 ;
        RECT 4.000 85.360 790.640 86.680 ;
        RECT 4.400 83.960 790.640 85.360 ;
        RECT 4.000 82.640 790.640 83.960 ;
        RECT 4.400 81.240 790.640 82.640 ;
        RECT 4.000 79.920 790.640 81.240 ;
        RECT 4.400 78.520 790.640 79.920 ;
        RECT 4.000 77.200 790.640 78.520 ;
        RECT 4.400 75.800 790.640 77.200 ;
        RECT 4.000 74.480 790.640 75.800 ;
        RECT 4.400 73.080 790.640 74.480 ;
        RECT 4.000 71.760 790.640 73.080 ;
        RECT 4.400 70.360 790.640 71.760 ;
        RECT 4.000 69.040 790.640 70.360 ;
        RECT 4.400 67.640 790.640 69.040 ;
        RECT 4.000 65.640 790.640 67.640 ;
        RECT 4.400 64.240 790.640 65.640 ;
        RECT 4.000 62.920 790.640 64.240 ;
        RECT 4.400 61.520 790.640 62.920 ;
        RECT 4.000 60.200 790.640 61.520 ;
        RECT 4.400 58.800 790.640 60.200 ;
        RECT 4.000 57.480 790.640 58.800 ;
        RECT 4.400 56.080 790.640 57.480 ;
        RECT 4.000 54.760 790.640 56.080 ;
        RECT 4.400 53.360 790.640 54.760 ;
        RECT 4.000 52.040 790.640 53.360 ;
        RECT 4.400 50.640 790.640 52.040 ;
        RECT 4.000 49.320 790.640 50.640 ;
        RECT 4.400 47.920 790.640 49.320 ;
        RECT 4.000 46.600 790.640 47.920 ;
        RECT 4.400 45.200 790.640 46.600 ;
        RECT 4.000 43.880 790.640 45.200 ;
        RECT 4.400 42.480 790.640 43.880 ;
        RECT 4.000 41.160 790.640 42.480 ;
        RECT 4.400 39.760 790.640 41.160 ;
        RECT 4.000 38.440 790.640 39.760 ;
        RECT 4.400 37.040 790.640 38.440 ;
        RECT 4.000 35.720 790.640 37.040 ;
        RECT 4.400 34.320 790.640 35.720 ;
        RECT 4.000 32.320 790.640 34.320 ;
        RECT 4.400 30.920 790.640 32.320 ;
        RECT 4.000 29.600 790.640 30.920 ;
        RECT 4.400 28.200 790.640 29.600 ;
        RECT 4.000 26.880 790.640 28.200 ;
        RECT 4.400 25.480 790.640 26.880 ;
        RECT 4.000 24.160 790.640 25.480 ;
        RECT 4.400 22.760 790.640 24.160 ;
        RECT 4.000 21.440 790.640 22.760 ;
        RECT 4.400 20.040 790.640 21.440 ;
        RECT 4.000 18.720 790.640 20.040 ;
        RECT 4.400 17.320 790.640 18.720 ;
        RECT 4.000 16.000 790.640 17.320 ;
        RECT 4.400 14.600 790.640 16.000 ;
        RECT 4.000 13.280 790.640 14.600 ;
        RECT 4.400 11.880 790.640 13.280 ;
        RECT 4.000 10.560 790.640 11.880 ;
        RECT 4.400 9.160 790.640 10.560 ;
        RECT 4.000 7.840 790.640 9.160 ;
        RECT 4.400 6.440 790.640 7.840 ;
        RECT 4.000 5.120 790.640 6.440 ;
        RECT 4.400 3.720 790.640 5.120 ;
        RECT 4.000 2.400 790.640 3.720 ;
        RECT 4.400 1.535 790.640 2.400 ;
      LAYER met4 ;
        RECT 11.335 288.960 759.625 299.705 ;
        RECT 11.335 134.135 20.640 288.960 ;
        RECT 23.040 134.135 97.440 288.960 ;
        RECT 99.840 134.135 174.240 288.960 ;
        RECT 176.640 134.135 251.040 288.960 ;
        RECT 253.440 134.135 327.840 288.960 ;
        RECT 330.240 134.135 404.640 288.960 ;
        RECT 407.040 134.135 481.440 288.960 ;
        RECT 483.840 134.135 558.240 288.960 ;
        RECT 560.640 134.135 635.040 288.960 ;
        RECT 637.440 134.135 711.840 288.960 ;
        RECT 714.240 134.135 759.625 288.960 ;
  END
END mkQF100Fabric
END LIBRARY

