magic
tech sky130A
magscale 1 2
timestamp 1647792197
<< obsli1 >>
rect 1104 2159 166980 167569
<< obsm1 >>
rect 14 2128 168070 168360
<< metal2 >>
rect 386 169453 442 170253
rect 1122 169453 1178 170253
rect 1950 169453 2006 170253
rect 2686 169453 2742 170253
rect 3514 169453 3570 170253
rect 4250 169453 4306 170253
rect 5078 169453 5134 170253
rect 5906 169453 5962 170253
rect 6642 169453 6698 170253
rect 7470 169453 7526 170253
rect 8206 169453 8262 170253
rect 9034 169453 9090 170253
rect 9770 169453 9826 170253
rect 10598 169453 10654 170253
rect 11426 169453 11482 170253
rect 12162 169453 12218 170253
rect 12990 169453 13046 170253
rect 13726 169453 13782 170253
rect 14554 169453 14610 170253
rect 15290 169453 15346 170253
rect 16118 169453 16174 170253
rect 16946 169453 17002 170253
rect 17682 169453 17738 170253
rect 18510 169453 18566 170253
rect 19246 169453 19302 170253
rect 20074 169453 20130 170253
rect 20902 169453 20958 170253
rect 21638 169453 21694 170253
rect 22466 169453 22522 170253
rect 23202 169453 23258 170253
rect 24030 169453 24086 170253
rect 24766 169453 24822 170253
rect 25594 169453 25650 170253
rect 26422 169453 26478 170253
rect 27158 169453 27214 170253
rect 27986 169453 28042 170253
rect 28722 169453 28778 170253
rect 29550 169453 29606 170253
rect 30286 169453 30342 170253
rect 31114 169453 31170 170253
rect 31942 169453 31998 170253
rect 32678 169453 32734 170253
rect 33506 169453 33562 170253
rect 34242 169453 34298 170253
rect 35070 169453 35126 170253
rect 35806 169453 35862 170253
rect 36634 169453 36690 170253
rect 37462 169453 37518 170253
rect 38198 169453 38254 170253
rect 39026 169453 39082 170253
rect 39762 169453 39818 170253
rect 40590 169453 40646 170253
rect 41418 169453 41474 170253
rect 42154 169453 42210 170253
rect 42982 169453 43038 170253
rect 43718 169453 43774 170253
rect 44546 169453 44602 170253
rect 45282 169453 45338 170253
rect 46110 169453 46166 170253
rect 46938 169453 46994 170253
rect 47674 169453 47730 170253
rect 48502 169453 48558 170253
rect 49238 169453 49294 170253
rect 50066 169453 50122 170253
rect 50802 169453 50858 170253
rect 51630 169453 51686 170253
rect 52458 169453 52514 170253
rect 53194 169453 53250 170253
rect 54022 169453 54078 170253
rect 54758 169453 54814 170253
rect 55586 169453 55642 170253
rect 56414 169453 56470 170253
rect 57150 169453 57206 170253
rect 57978 169453 58034 170253
rect 58714 169453 58770 170253
rect 59542 169453 59598 170253
rect 60278 169453 60334 170253
rect 61106 169453 61162 170253
rect 61934 169453 61990 170253
rect 62670 169453 62726 170253
rect 63498 169453 63554 170253
rect 64234 169453 64290 170253
rect 65062 169453 65118 170253
rect 65798 169453 65854 170253
rect 66626 169453 66682 170253
rect 67454 169453 67510 170253
rect 68190 169453 68246 170253
rect 69018 169453 69074 170253
rect 69754 169453 69810 170253
rect 70582 169453 70638 170253
rect 71318 169453 71374 170253
rect 72146 169453 72202 170253
rect 72974 169453 73030 170253
rect 73710 169453 73766 170253
rect 74538 169453 74594 170253
rect 75274 169453 75330 170253
rect 76102 169453 76158 170253
rect 76930 169453 76986 170253
rect 77666 169453 77722 170253
rect 78494 169453 78550 170253
rect 79230 169453 79286 170253
rect 80058 169453 80114 170253
rect 80794 169453 80850 170253
rect 81622 169453 81678 170253
rect 82450 169453 82506 170253
rect 83186 169453 83242 170253
rect 84014 169453 84070 170253
rect 84750 169453 84806 170253
rect 85578 169453 85634 170253
rect 86314 169453 86370 170253
rect 87142 169453 87198 170253
rect 87970 169453 88026 170253
rect 88706 169453 88762 170253
rect 89534 169453 89590 170253
rect 90270 169453 90326 170253
rect 91098 169453 91154 170253
rect 91834 169453 91890 170253
rect 92662 169453 92718 170253
rect 93490 169453 93546 170253
rect 94226 169453 94282 170253
rect 95054 169453 95110 170253
rect 95790 169453 95846 170253
rect 96618 169453 96674 170253
rect 97446 169453 97502 170253
rect 98182 169453 98238 170253
rect 99010 169453 99066 170253
rect 99746 169453 99802 170253
rect 100574 169453 100630 170253
rect 101310 169453 101366 170253
rect 102138 169453 102194 170253
rect 102966 169453 103022 170253
rect 103702 169453 103758 170253
rect 104530 169453 104586 170253
rect 105266 169453 105322 170253
rect 106094 169453 106150 170253
rect 106830 169453 106886 170253
rect 107658 169453 107714 170253
rect 108486 169453 108542 170253
rect 109222 169453 109278 170253
rect 110050 169453 110106 170253
rect 110786 169453 110842 170253
rect 111614 169453 111670 170253
rect 112442 169453 112498 170253
rect 113178 169453 113234 170253
rect 114006 169453 114062 170253
rect 114742 169453 114798 170253
rect 115570 169453 115626 170253
rect 116306 169453 116362 170253
rect 117134 169453 117190 170253
rect 117962 169453 118018 170253
rect 118698 169453 118754 170253
rect 119526 169453 119582 170253
rect 120262 169453 120318 170253
rect 121090 169453 121146 170253
rect 121826 169453 121882 170253
rect 122654 169453 122710 170253
rect 123482 169453 123538 170253
rect 124218 169453 124274 170253
rect 125046 169453 125102 170253
rect 125782 169453 125838 170253
rect 126610 169453 126666 170253
rect 127346 169453 127402 170253
rect 128174 169453 128230 170253
rect 129002 169453 129058 170253
rect 129738 169453 129794 170253
rect 130566 169453 130622 170253
rect 131302 169453 131358 170253
rect 132130 169453 132186 170253
rect 132958 169453 133014 170253
rect 133694 169453 133750 170253
rect 134522 169453 134578 170253
rect 135258 169453 135314 170253
rect 136086 169453 136142 170253
rect 136822 169453 136878 170253
rect 137650 169453 137706 170253
rect 138478 169453 138534 170253
rect 139214 169453 139270 170253
rect 140042 169453 140098 170253
rect 140778 169453 140834 170253
rect 141606 169453 141662 170253
rect 142342 169453 142398 170253
rect 143170 169453 143226 170253
rect 143998 169453 144054 170253
rect 144734 169453 144790 170253
rect 145562 169453 145618 170253
rect 146298 169453 146354 170253
rect 147126 169453 147182 170253
rect 147862 169453 147918 170253
rect 148690 169453 148746 170253
rect 149518 169453 149574 170253
rect 150254 169453 150310 170253
rect 151082 169453 151138 170253
rect 151818 169453 151874 170253
rect 152646 169453 152702 170253
rect 153474 169453 153530 170253
rect 154210 169453 154266 170253
rect 155038 169453 155094 170253
rect 155774 169453 155830 170253
rect 156602 169453 156658 170253
rect 157338 169453 157394 170253
rect 158166 169453 158222 170253
rect 158994 169453 159050 170253
rect 159730 169453 159786 170253
rect 160558 169453 160614 170253
rect 161294 169453 161350 170253
rect 162122 169453 162178 170253
rect 162858 169453 162914 170253
rect 163686 169453 163742 170253
rect 164514 169453 164570 170253
rect 165250 169453 165306 170253
rect 166078 169453 166134 170253
rect 166814 169453 166870 170253
rect 167642 169453 167698 170253
rect 9310 0 9366 800
rect 27986 0 28042 800
rect 46662 0 46718 800
rect 65338 0 65394 800
rect 84014 0 84070 800
rect 102690 0 102746 800
rect 121366 0 121422 800
rect 140042 0 140098 800
rect 158718 0 158774 800
<< obsm2 >>
rect 20 169397 330 169538
rect 498 169397 1066 169538
rect 1234 169397 1894 169538
rect 2062 169397 2630 169538
rect 2798 169397 3458 169538
rect 3626 169397 4194 169538
rect 4362 169397 5022 169538
rect 5190 169397 5850 169538
rect 6018 169397 6586 169538
rect 6754 169397 7414 169538
rect 7582 169397 8150 169538
rect 8318 169397 8978 169538
rect 9146 169397 9714 169538
rect 9882 169397 10542 169538
rect 10710 169397 11370 169538
rect 11538 169397 12106 169538
rect 12274 169397 12934 169538
rect 13102 169397 13670 169538
rect 13838 169397 14498 169538
rect 14666 169397 15234 169538
rect 15402 169397 16062 169538
rect 16230 169397 16890 169538
rect 17058 169397 17626 169538
rect 17794 169397 18454 169538
rect 18622 169397 19190 169538
rect 19358 169397 20018 169538
rect 20186 169397 20846 169538
rect 21014 169397 21582 169538
rect 21750 169397 22410 169538
rect 22578 169397 23146 169538
rect 23314 169397 23974 169538
rect 24142 169397 24710 169538
rect 24878 169397 25538 169538
rect 25706 169397 26366 169538
rect 26534 169397 27102 169538
rect 27270 169397 27930 169538
rect 28098 169397 28666 169538
rect 28834 169397 29494 169538
rect 29662 169397 30230 169538
rect 30398 169397 31058 169538
rect 31226 169397 31886 169538
rect 32054 169397 32622 169538
rect 32790 169397 33450 169538
rect 33618 169397 34186 169538
rect 34354 169397 35014 169538
rect 35182 169397 35750 169538
rect 35918 169397 36578 169538
rect 36746 169397 37406 169538
rect 37574 169397 38142 169538
rect 38310 169397 38970 169538
rect 39138 169397 39706 169538
rect 39874 169397 40534 169538
rect 40702 169397 41362 169538
rect 41530 169397 42098 169538
rect 42266 169397 42926 169538
rect 43094 169397 43662 169538
rect 43830 169397 44490 169538
rect 44658 169397 45226 169538
rect 45394 169397 46054 169538
rect 46222 169397 46882 169538
rect 47050 169397 47618 169538
rect 47786 169397 48446 169538
rect 48614 169397 49182 169538
rect 49350 169397 50010 169538
rect 50178 169397 50746 169538
rect 50914 169397 51574 169538
rect 51742 169397 52402 169538
rect 52570 169397 53138 169538
rect 53306 169397 53966 169538
rect 54134 169397 54702 169538
rect 54870 169397 55530 169538
rect 55698 169397 56358 169538
rect 56526 169397 57094 169538
rect 57262 169397 57922 169538
rect 58090 169397 58658 169538
rect 58826 169397 59486 169538
rect 59654 169397 60222 169538
rect 60390 169397 61050 169538
rect 61218 169397 61878 169538
rect 62046 169397 62614 169538
rect 62782 169397 63442 169538
rect 63610 169397 64178 169538
rect 64346 169397 65006 169538
rect 65174 169397 65742 169538
rect 65910 169397 66570 169538
rect 66738 169397 67398 169538
rect 67566 169397 68134 169538
rect 68302 169397 68962 169538
rect 69130 169397 69698 169538
rect 69866 169397 70526 169538
rect 70694 169397 71262 169538
rect 71430 169397 72090 169538
rect 72258 169397 72918 169538
rect 73086 169397 73654 169538
rect 73822 169397 74482 169538
rect 74650 169397 75218 169538
rect 75386 169397 76046 169538
rect 76214 169397 76874 169538
rect 77042 169397 77610 169538
rect 77778 169397 78438 169538
rect 78606 169397 79174 169538
rect 79342 169397 80002 169538
rect 80170 169397 80738 169538
rect 80906 169397 81566 169538
rect 81734 169397 82394 169538
rect 82562 169397 83130 169538
rect 83298 169397 83958 169538
rect 84126 169397 84694 169538
rect 84862 169397 85522 169538
rect 85690 169397 86258 169538
rect 86426 169397 87086 169538
rect 87254 169397 87914 169538
rect 88082 169397 88650 169538
rect 88818 169397 89478 169538
rect 89646 169397 90214 169538
rect 90382 169397 91042 169538
rect 91210 169397 91778 169538
rect 91946 169397 92606 169538
rect 92774 169397 93434 169538
rect 93602 169397 94170 169538
rect 94338 169397 94998 169538
rect 95166 169397 95734 169538
rect 95902 169397 96562 169538
rect 96730 169397 97390 169538
rect 97558 169397 98126 169538
rect 98294 169397 98954 169538
rect 99122 169397 99690 169538
rect 99858 169397 100518 169538
rect 100686 169397 101254 169538
rect 101422 169397 102082 169538
rect 102250 169397 102910 169538
rect 103078 169397 103646 169538
rect 103814 169397 104474 169538
rect 104642 169397 105210 169538
rect 105378 169397 106038 169538
rect 106206 169397 106774 169538
rect 106942 169397 107602 169538
rect 107770 169397 108430 169538
rect 108598 169397 109166 169538
rect 109334 169397 109994 169538
rect 110162 169397 110730 169538
rect 110898 169397 111558 169538
rect 111726 169397 112386 169538
rect 112554 169397 113122 169538
rect 113290 169397 113950 169538
rect 114118 169397 114686 169538
rect 114854 169397 115514 169538
rect 115682 169397 116250 169538
rect 116418 169397 117078 169538
rect 117246 169397 117906 169538
rect 118074 169397 118642 169538
rect 118810 169397 119470 169538
rect 119638 169397 120206 169538
rect 120374 169397 121034 169538
rect 121202 169397 121770 169538
rect 121938 169397 122598 169538
rect 122766 169397 123426 169538
rect 123594 169397 124162 169538
rect 124330 169397 124990 169538
rect 125158 169397 125726 169538
rect 125894 169397 126554 169538
rect 126722 169397 127290 169538
rect 127458 169397 128118 169538
rect 128286 169397 128946 169538
rect 129114 169397 129682 169538
rect 129850 169397 130510 169538
rect 130678 169397 131246 169538
rect 131414 169397 132074 169538
rect 132242 169397 132902 169538
rect 133070 169397 133638 169538
rect 133806 169397 134466 169538
rect 134634 169397 135202 169538
rect 135370 169397 136030 169538
rect 136198 169397 136766 169538
rect 136934 169397 137594 169538
rect 137762 169397 138422 169538
rect 138590 169397 139158 169538
rect 139326 169397 139986 169538
rect 140154 169397 140722 169538
rect 140890 169397 141550 169538
rect 141718 169397 142286 169538
rect 142454 169397 143114 169538
rect 143282 169397 143942 169538
rect 144110 169397 144678 169538
rect 144846 169397 145506 169538
rect 145674 169397 146242 169538
rect 146410 169397 147070 169538
rect 147238 169397 147806 169538
rect 147974 169397 148634 169538
rect 148802 169397 149462 169538
rect 149630 169397 150198 169538
rect 150366 169397 151026 169538
rect 151194 169397 151762 169538
rect 151930 169397 152590 169538
rect 152758 169397 153418 169538
rect 153586 169397 154154 169538
rect 154322 169397 154982 169538
rect 155150 169397 155718 169538
rect 155886 169397 156546 169538
rect 156714 169397 157282 169538
rect 157450 169397 158110 169538
rect 158278 169397 158938 169538
rect 159106 169397 159674 169538
rect 159842 169397 160502 169538
rect 160670 169397 161238 169538
rect 161406 169397 162066 169538
rect 162234 169397 162802 169538
rect 162970 169397 163630 169538
rect 163798 169397 164458 169538
rect 164626 169397 165194 169538
rect 165362 169397 166022 169538
rect 166190 169397 166758 169538
rect 166926 169397 167586 169538
rect 167754 169397 168064 169538
rect 20 856 168064 169397
rect 20 711 9254 856
rect 9422 711 27930 856
rect 28098 711 46606 856
rect 46774 711 65282 856
rect 65450 711 83958 856
rect 84126 711 102634 856
rect 102802 711 121310 856
rect 121478 711 139986 856
rect 140154 711 158662 856
rect 158830 711 168064 856
<< metal3 >>
rect 167309 169328 168109 169448
rect 167309 167832 168109 167952
rect 167309 166336 168109 166456
rect 167309 164840 168109 164960
rect 167309 163344 168109 163464
rect 167309 161848 168109 161968
rect 0 161576 800 161696
rect 167309 160352 168109 160472
rect 167309 158856 168109 158976
rect 167309 157360 168109 157480
rect 167309 155864 168109 155984
rect 167309 154368 168109 154488
rect 167309 152872 168109 152992
rect 167309 151240 168109 151360
rect 167309 149744 168109 149864
rect 167309 148248 168109 148368
rect 167309 146752 168109 146872
rect 167309 145256 168109 145376
rect 0 144576 800 144696
rect 167309 143760 168109 143880
rect 167309 142264 168109 142384
rect 167309 140768 168109 140888
rect 167309 139272 168109 139392
rect 167309 137776 168109 137896
rect 167309 136280 168109 136400
rect 167309 134784 168109 134904
rect 167309 133288 168109 133408
rect 167309 131656 168109 131776
rect 167309 130160 168109 130280
rect 167309 128664 168109 128784
rect 0 127576 800 127696
rect 167309 127168 168109 127288
rect 167309 125672 168109 125792
rect 167309 124176 168109 124296
rect 167309 122680 168109 122800
rect 167309 121184 168109 121304
rect 167309 119688 168109 119808
rect 167309 118192 168109 118312
rect 167309 116696 168109 116816
rect 167309 115200 168109 115320
rect 167309 113568 168109 113688
rect 167309 112072 168109 112192
rect 0 110576 800 110696
rect 167309 110576 168109 110696
rect 167309 109080 168109 109200
rect 167309 107584 168109 107704
rect 167309 106088 168109 106208
rect 167309 104592 168109 104712
rect 167309 103096 168109 103216
rect 167309 101600 168109 101720
rect 167309 100104 168109 100224
rect 167309 98608 168109 98728
rect 167309 97112 168109 97232
rect 167309 95616 168109 95736
rect 167309 93984 168109 94104
rect 0 93576 800 93696
rect 167309 92488 168109 92608
rect 167309 90992 168109 91112
rect 167309 89496 168109 89616
rect 167309 88000 168109 88120
rect 167309 86504 168109 86624
rect 167309 85008 168109 85128
rect 167309 83512 168109 83632
rect 167309 82016 168109 82136
rect 167309 80520 168109 80640
rect 167309 79024 168109 79144
rect 167309 77528 168109 77648
rect 0 76440 800 76560
rect 167309 75896 168109 76016
rect 167309 74400 168109 74520
rect 167309 72904 168109 73024
rect 167309 71408 168109 71528
rect 167309 69912 168109 70032
rect 167309 68416 168109 68536
rect 167309 66920 168109 67040
rect 167309 65424 168109 65544
rect 167309 63928 168109 64048
rect 167309 62432 168109 62552
rect 167309 60936 168109 61056
rect 0 59440 800 59560
rect 167309 59440 168109 59560
rect 167309 57944 168109 58064
rect 167309 56312 168109 56432
rect 167309 54816 168109 54936
rect 167309 53320 168109 53440
rect 167309 51824 168109 51944
rect 167309 50328 168109 50448
rect 167309 48832 168109 48952
rect 167309 47336 168109 47456
rect 167309 45840 168109 45960
rect 167309 44344 168109 44464
rect 167309 42848 168109 42968
rect 0 42440 800 42560
rect 167309 41352 168109 41472
rect 167309 39856 168109 39976
rect 167309 38224 168109 38344
rect 167309 36728 168109 36848
rect 167309 35232 168109 35352
rect 167309 33736 168109 33856
rect 167309 32240 168109 32360
rect 167309 30744 168109 30864
rect 167309 29248 168109 29368
rect 167309 27752 168109 27872
rect 167309 26256 168109 26376
rect 0 25440 800 25560
rect 167309 24760 168109 24880
rect 167309 23264 168109 23384
rect 167309 21768 168109 21888
rect 167309 20272 168109 20392
rect 167309 18640 168109 18760
rect 167309 17144 168109 17264
rect 167309 15648 168109 15768
rect 167309 14152 168109 14272
rect 167309 12656 168109 12776
rect 167309 11160 168109 11280
rect 167309 9664 168109 9784
rect 0 8440 800 8560
rect 167309 8168 168109 8288
rect 167309 6672 168109 6792
rect 167309 5176 168109 5296
rect 167309 3680 168109 3800
rect 167309 2184 168109 2304
rect 167309 688 168109 808
<< obsm3 >>
rect 800 169248 167229 169421
rect 800 168032 167378 169248
rect 800 167752 167229 168032
rect 800 166536 167378 167752
rect 800 166256 167229 166536
rect 800 165040 167378 166256
rect 800 164760 167229 165040
rect 800 163544 167378 164760
rect 800 163264 167229 163544
rect 800 162048 167378 163264
rect 800 161776 167229 162048
rect 880 161768 167229 161776
rect 880 161496 167378 161768
rect 800 160552 167378 161496
rect 800 160272 167229 160552
rect 800 159056 167378 160272
rect 800 158776 167229 159056
rect 800 157560 167378 158776
rect 800 157280 167229 157560
rect 800 156064 167378 157280
rect 800 155784 167229 156064
rect 800 154568 167378 155784
rect 800 154288 167229 154568
rect 800 153072 167378 154288
rect 800 152792 167229 153072
rect 800 151440 167378 152792
rect 800 151160 167229 151440
rect 800 149944 167378 151160
rect 800 149664 167229 149944
rect 800 148448 167378 149664
rect 800 148168 167229 148448
rect 800 146952 167378 148168
rect 800 146672 167229 146952
rect 800 145456 167378 146672
rect 800 145176 167229 145456
rect 800 144776 167378 145176
rect 880 144496 167378 144776
rect 800 143960 167378 144496
rect 800 143680 167229 143960
rect 800 142464 167378 143680
rect 800 142184 167229 142464
rect 800 140968 167378 142184
rect 800 140688 167229 140968
rect 800 139472 167378 140688
rect 800 139192 167229 139472
rect 800 137976 167378 139192
rect 800 137696 167229 137976
rect 800 136480 167378 137696
rect 800 136200 167229 136480
rect 800 134984 167378 136200
rect 800 134704 167229 134984
rect 800 133488 167378 134704
rect 800 133208 167229 133488
rect 800 131856 167378 133208
rect 800 131576 167229 131856
rect 800 130360 167378 131576
rect 800 130080 167229 130360
rect 800 128864 167378 130080
rect 800 128584 167229 128864
rect 800 127776 167378 128584
rect 880 127496 167378 127776
rect 800 127368 167378 127496
rect 800 127088 167229 127368
rect 800 125872 167378 127088
rect 800 125592 167229 125872
rect 800 124376 167378 125592
rect 800 124096 167229 124376
rect 800 122880 167378 124096
rect 800 122600 167229 122880
rect 800 121384 167378 122600
rect 800 121104 167229 121384
rect 800 119888 167378 121104
rect 800 119608 167229 119888
rect 800 118392 167378 119608
rect 800 118112 167229 118392
rect 800 116896 167378 118112
rect 800 116616 167229 116896
rect 800 115400 167378 116616
rect 800 115120 167229 115400
rect 800 113768 167378 115120
rect 800 113488 167229 113768
rect 800 112272 167378 113488
rect 800 111992 167229 112272
rect 800 110776 167378 111992
rect 880 110496 167229 110776
rect 800 109280 167378 110496
rect 800 109000 167229 109280
rect 800 107784 167378 109000
rect 800 107504 167229 107784
rect 800 106288 167378 107504
rect 800 106008 167229 106288
rect 800 104792 167378 106008
rect 800 104512 167229 104792
rect 800 103296 167378 104512
rect 800 103016 167229 103296
rect 800 101800 167378 103016
rect 800 101520 167229 101800
rect 800 100304 167378 101520
rect 800 100024 167229 100304
rect 800 98808 167378 100024
rect 800 98528 167229 98808
rect 800 97312 167378 98528
rect 800 97032 167229 97312
rect 800 95816 167378 97032
rect 800 95536 167229 95816
rect 800 94184 167378 95536
rect 800 93904 167229 94184
rect 800 93776 167378 93904
rect 880 93496 167378 93776
rect 800 92688 167378 93496
rect 800 92408 167229 92688
rect 800 91192 167378 92408
rect 800 90912 167229 91192
rect 800 89696 167378 90912
rect 800 89416 167229 89696
rect 800 88200 167378 89416
rect 800 87920 167229 88200
rect 800 86704 167378 87920
rect 800 86424 167229 86704
rect 800 85208 167378 86424
rect 800 84928 167229 85208
rect 800 83712 167378 84928
rect 800 83432 167229 83712
rect 800 82216 167378 83432
rect 800 81936 167229 82216
rect 800 80720 167378 81936
rect 800 80440 167229 80720
rect 800 79224 167378 80440
rect 800 78944 167229 79224
rect 800 77728 167378 78944
rect 800 77448 167229 77728
rect 800 76640 167378 77448
rect 880 76360 167378 76640
rect 800 76096 167378 76360
rect 800 75816 167229 76096
rect 800 74600 167378 75816
rect 800 74320 167229 74600
rect 800 73104 167378 74320
rect 800 72824 167229 73104
rect 800 71608 167378 72824
rect 800 71328 167229 71608
rect 800 70112 167378 71328
rect 800 69832 167229 70112
rect 800 68616 167378 69832
rect 800 68336 167229 68616
rect 800 67120 167378 68336
rect 800 66840 167229 67120
rect 800 65624 167378 66840
rect 800 65344 167229 65624
rect 800 64128 167378 65344
rect 800 63848 167229 64128
rect 800 62632 167378 63848
rect 800 62352 167229 62632
rect 800 61136 167378 62352
rect 800 60856 167229 61136
rect 800 59640 167378 60856
rect 880 59360 167229 59640
rect 800 58144 167378 59360
rect 800 57864 167229 58144
rect 800 56512 167378 57864
rect 800 56232 167229 56512
rect 800 55016 167378 56232
rect 800 54736 167229 55016
rect 800 53520 167378 54736
rect 800 53240 167229 53520
rect 800 52024 167378 53240
rect 800 51744 167229 52024
rect 800 50528 167378 51744
rect 800 50248 167229 50528
rect 800 49032 167378 50248
rect 800 48752 167229 49032
rect 800 47536 167378 48752
rect 800 47256 167229 47536
rect 800 46040 167378 47256
rect 800 45760 167229 46040
rect 800 44544 167378 45760
rect 800 44264 167229 44544
rect 800 43048 167378 44264
rect 800 42768 167229 43048
rect 800 42640 167378 42768
rect 880 42360 167378 42640
rect 800 41552 167378 42360
rect 800 41272 167229 41552
rect 800 40056 167378 41272
rect 800 39776 167229 40056
rect 800 38424 167378 39776
rect 800 38144 167229 38424
rect 800 36928 167378 38144
rect 800 36648 167229 36928
rect 800 35432 167378 36648
rect 800 35152 167229 35432
rect 800 33936 167378 35152
rect 800 33656 167229 33936
rect 800 32440 167378 33656
rect 800 32160 167229 32440
rect 800 30944 167378 32160
rect 800 30664 167229 30944
rect 800 29448 167378 30664
rect 800 29168 167229 29448
rect 800 27952 167378 29168
rect 800 27672 167229 27952
rect 800 26456 167378 27672
rect 800 26176 167229 26456
rect 800 25640 167378 26176
rect 880 25360 167378 25640
rect 800 24960 167378 25360
rect 800 24680 167229 24960
rect 800 23464 167378 24680
rect 800 23184 167229 23464
rect 800 21968 167378 23184
rect 800 21688 167229 21968
rect 800 20472 167378 21688
rect 800 20192 167229 20472
rect 800 18840 167378 20192
rect 800 18560 167229 18840
rect 800 17344 167378 18560
rect 800 17064 167229 17344
rect 800 15848 167378 17064
rect 800 15568 167229 15848
rect 800 14352 167378 15568
rect 800 14072 167229 14352
rect 800 12856 167378 14072
rect 800 12576 167229 12856
rect 800 11360 167378 12576
rect 800 11080 167229 11360
rect 800 9864 167378 11080
rect 800 9584 167229 9864
rect 800 8640 167378 9584
rect 880 8368 167378 8640
rect 880 8360 167229 8368
rect 800 8088 167229 8360
rect 800 6872 167378 8088
rect 800 6592 167229 6872
rect 800 5376 167378 6592
rect 800 5096 167229 5376
rect 800 3880 167378 5096
rect 800 3600 167229 3880
rect 800 2384 167378 3600
rect 800 2104 167229 2384
rect 800 888 167378 2104
rect 800 715 167229 888
<< metal4 >>
rect 4208 2128 4528 167600
rect 19568 2128 19888 167600
rect 34928 2128 35248 167600
rect 50288 2128 50608 167600
rect 65648 2128 65968 167600
rect 81008 2128 81328 167600
rect 96368 2128 96688 167600
rect 111728 2128 112048 167600
rect 127088 2128 127408 167600
rect 142448 2128 142768 167600
rect 157808 2128 158128 167600
<< obsm4 >>
rect 4659 3299 19488 165749
rect 19968 3299 34848 165749
rect 35328 3299 50208 165749
rect 50688 3299 65568 165749
rect 66048 3299 80928 165749
rect 81408 3299 96288 165749
rect 96768 3299 111648 165749
rect 112128 3299 127008 165749
rect 127488 3299 142368 165749
rect 142848 3299 157728 165749
rect 158208 3299 165541 165749
<< labels >>
rlabel metal2 s 27986 0 28042 800 6 CLK
port 1 nsew signal input
rlabel metal2 s 386 169453 442 170253 6 EN_dmem_client_request_get
port 2 nsew signal input
rlabel metal2 s 1122 169453 1178 170253 6 EN_dmem_client_response_put
port 3 nsew signal input
rlabel metal2 s 107658 169453 107714 170253 6 EN_imem_client_request_get
port 4 nsew signal input
rlabel metal2 s 108486 169453 108542 170253 6 EN_imem_client_response_put
port 5 nsew signal input
rlabel metal2 s 1950 169453 2006 170253 6 RDY_dmem_client_request_get
port 6 nsew signal output
rlabel metal2 s 2686 169453 2742 170253 6 RDY_dmem_client_response_put
port 7 nsew signal output
rlabel metal2 s 109222 169453 109278 170253 6 RDY_imem_client_request_get
port 8 nsew signal output
rlabel metal2 s 110050 169453 110106 170253 6 RDY_imem_client_response_put
port 9 nsew signal output
rlabel metal2 s 46662 0 46718 800 6 RDY_readPC
port 10 nsew signal output
rlabel metal2 s 9310 0 9366 800 6 RST_N
port 11 nsew signal input
rlabel metal2 s 3514 169453 3570 170253 6 dmem_client_request_get[0]
port 12 nsew signal output
rlabel metal2 s 19246 169453 19302 170253 6 dmem_client_request_get[10]
port 13 nsew signal output
rlabel metal2 s 20902 169453 20958 170253 6 dmem_client_request_get[11]
port 14 nsew signal output
rlabel metal2 s 22466 169453 22522 170253 6 dmem_client_request_get[12]
port 15 nsew signal output
rlabel metal2 s 24030 169453 24086 170253 6 dmem_client_request_get[13]
port 16 nsew signal output
rlabel metal2 s 25594 169453 25650 170253 6 dmem_client_request_get[14]
port 17 nsew signal output
rlabel metal2 s 27158 169453 27214 170253 6 dmem_client_request_get[15]
port 18 nsew signal output
rlabel metal2 s 28722 169453 28778 170253 6 dmem_client_request_get[16]
port 19 nsew signal output
rlabel metal2 s 30286 169453 30342 170253 6 dmem_client_request_get[17]
port 20 nsew signal output
rlabel metal2 s 31942 169453 31998 170253 6 dmem_client_request_get[18]
port 21 nsew signal output
rlabel metal2 s 33506 169453 33562 170253 6 dmem_client_request_get[19]
port 22 nsew signal output
rlabel metal2 s 5078 169453 5134 170253 6 dmem_client_request_get[1]
port 23 nsew signal output
rlabel metal2 s 35070 169453 35126 170253 6 dmem_client_request_get[20]
port 24 nsew signal output
rlabel metal2 s 36634 169453 36690 170253 6 dmem_client_request_get[21]
port 25 nsew signal output
rlabel metal2 s 38198 169453 38254 170253 6 dmem_client_request_get[22]
port 26 nsew signal output
rlabel metal2 s 39762 169453 39818 170253 6 dmem_client_request_get[23]
port 27 nsew signal output
rlabel metal2 s 41418 169453 41474 170253 6 dmem_client_request_get[24]
port 28 nsew signal output
rlabel metal2 s 42982 169453 43038 170253 6 dmem_client_request_get[25]
port 29 nsew signal output
rlabel metal2 s 44546 169453 44602 170253 6 dmem_client_request_get[26]
port 30 nsew signal output
rlabel metal2 s 46110 169453 46166 170253 6 dmem_client_request_get[27]
port 31 nsew signal output
rlabel metal2 s 47674 169453 47730 170253 6 dmem_client_request_get[28]
port 32 nsew signal output
rlabel metal2 s 49238 169453 49294 170253 6 dmem_client_request_get[29]
port 33 nsew signal output
rlabel metal2 s 6642 169453 6698 170253 6 dmem_client_request_get[2]
port 34 nsew signal output
rlabel metal2 s 50802 169453 50858 170253 6 dmem_client_request_get[30]
port 35 nsew signal output
rlabel metal2 s 52458 169453 52514 170253 6 dmem_client_request_get[31]
port 36 nsew signal output
rlabel metal2 s 54022 169453 54078 170253 6 dmem_client_request_get[32]
port 37 nsew signal output
rlabel metal2 s 54758 169453 54814 170253 6 dmem_client_request_get[33]
port 38 nsew signal output
rlabel metal2 s 55586 169453 55642 170253 6 dmem_client_request_get[34]
port 39 nsew signal output
rlabel metal2 s 56414 169453 56470 170253 6 dmem_client_request_get[35]
port 40 nsew signal output
rlabel metal2 s 57150 169453 57206 170253 6 dmem_client_request_get[36]
port 41 nsew signal output
rlabel metal2 s 57978 169453 58034 170253 6 dmem_client_request_get[37]
port 42 nsew signal output
rlabel metal2 s 58714 169453 58770 170253 6 dmem_client_request_get[38]
port 43 nsew signal output
rlabel metal2 s 59542 169453 59598 170253 6 dmem_client_request_get[39]
port 44 nsew signal output
rlabel metal2 s 8206 169453 8262 170253 6 dmem_client_request_get[3]
port 45 nsew signal output
rlabel metal2 s 60278 169453 60334 170253 6 dmem_client_request_get[40]
port 46 nsew signal output
rlabel metal2 s 61106 169453 61162 170253 6 dmem_client_request_get[41]
port 47 nsew signal output
rlabel metal2 s 61934 169453 61990 170253 6 dmem_client_request_get[42]
port 48 nsew signal output
rlabel metal2 s 62670 169453 62726 170253 6 dmem_client_request_get[43]
port 49 nsew signal output
rlabel metal2 s 63498 169453 63554 170253 6 dmem_client_request_get[44]
port 50 nsew signal output
rlabel metal2 s 64234 169453 64290 170253 6 dmem_client_request_get[45]
port 51 nsew signal output
rlabel metal2 s 65062 169453 65118 170253 6 dmem_client_request_get[46]
port 52 nsew signal output
rlabel metal2 s 65798 169453 65854 170253 6 dmem_client_request_get[47]
port 53 nsew signal output
rlabel metal2 s 66626 169453 66682 170253 6 dmem_client_request_get[48]
port 54 nsew signal output
rlabel metal2 s 67454 169453 67510 170253 6 dmem_client_request_get[49]
port 55 nsew signal output
rlabel metal2 s 9770 169453 9826 170253 6 dmem_client_request_get[4]
port 56 nsew signal output
rlabel metal2 s 68190 169453 68246 170253 6 dmem_client_request_get[50]
port 57 nsew signal output
rlabel metal2 s 69018 169453 69074 170253 6 dmem_client_request_get[51]
port 58 nsew signal output
rlabel metal2 s 69754 169453 69810 170253 6 dmem_client_request_get[52]
port 59 nsew signal output
rlabel metal2 s 70582 169453 70638 170253 6 dmem_client_request_get[53]
port 60 nsew signal output
rlabel metal2 s 71318 169453 71374 170253 6 dmem_client_request_get[54]
port 61 nsew signal output
rlabel metal2 s 72146 169453 72202 170253 6 dmem_client_request_get[55]
port 62 nsew signal output
rlabel metal2 s 72974 169453 73030 170253 6 dmem_client_request_get[56]
port 63 nsew signal output
rlabel metal2 s 73710 169453 73766 170253 6 dmem_client_request_get[57]
port 64 nsew signal output
rlabel metal2 s 74538 169453 74594 170253 6 dmem_client_request_get[58]
port 65 nsew signal output
rlabel metal2 s 75274 169453 75330 170253 6 dmem_client_request_get[59]
port 66 nsew signal output
rlabel metal2 s 11426 169453 11482 170253 6 dmem_client_request_get[5]
port 67 nsew signal output
rlabel metal2 s 76102 169453 76158 170253 6 dmem_client_request_get[60]
port 68 nsew signal output
rlabel metal2 s 76930 169453 76986 170253 6 dmem_client_request_get[61]
port 69 nsew signal output
rlabel metal2 s 77666 169453 77722 170253 6 dmem_client_request_get[62]
port 70 nsew signal output
rlabel metal2 s 78494 169453 78550 170253 6 dmem_client_request_get[63]
port 71 nsew signal output
rlabel metal2 s 79230 169453 79286 170253 6 dmem_client_request_get[64]
port 72 nsew signal output
rlabel metal2 s 80058 169453 80114 170253 6 dmem_client_request_get[65]
port 73 nsew signal output
rlabel metal2 s 80794 169453 80850 170253 6 dmem_client_request_get[66]
port 74 nsew signal output
rlabel metal2 s 81622 169453 81678 170253 6 dmem_client_request_get[67]
port 75 nsew signal output
rlabel metal2 s 82450 169453 82506 170253 6 dmem_client_request_get[68]
port 76 nsew signal output
rlabel metal2 s 83186 169453 83242 170253 6 dmem_client_request_get[69]
port 77 nsew signal output
rlabel metal2 s 12990 169453 13046 170253 6 dmem_client_request_get[6]
port 78 nsew signal output
rlabel metal2 s 84014 169453 84070 170253 6 dmem_client_request_get[70]
port 79 nsew signal output
rlabel metal2 s 84750 169453 84806 170253 6 dmem_client_request_get[71]
port 80 nsew signal output
rlabel metal2 s 85578 169453 85634 170253 6 dmem_client_request_get[72]
port 81 nsew signal output
rlabel metal2 s 86314 169453 86370 170253 6 dmem_client_request_get[73]
port 82 nsew signal output
rlabel metal2 s 87142 169453 87198 170253 6 dmem_client_request_get[74]
port 83 nsew signal output
rlabel metal2 s 87970 169453 88026 170253 6 dmem_client_request_get[75]
port 84 nsew signal output
rlabel metal2 s 88706 169453 88762 170253 6 dmem_client_request_get[76]
port 85 nsew signal output
rlabel metal2 s 89534 169453 89590 170253 6 dmem_client_request_get[77]
port 86 nsew signal output
rlabel metal2 s 90270 169453 90326 170253 6 dmem_client_request_get[78]
port 87 nsew signal output
rlabel metal2 s 91098 169453 91154 170253 6 dmem_client_request_get[79]
port 88 nsew signal output
rlabel metal2 s 14554 169453 14610 170253 6 dmem_client_request_get[7]
port 89 nsew signal output
rlabel metal2 s 91834 169453 91890 170253 6 dmem_client_request_get[80]
port 90 nsew signal output
rlabel metal2 s 92662 169453 92718 170253 6 dmem_client_request_get[81]
port 91 nsew signal output
rlabel metal2 s 93490 169453 93546 170253 6 dmem_client_request_get[82]
port 92 nsew signal output
rlabel metal2 s 94226 169453 94282 170253 6 dmem_client_request_get[83]
port 93 nsew signal output
rlabel metal2 s 95054 169453 95110 170253 6 dmem_client_request_get[84]
port 94 nsew signal output
rlabel metal2 s 95790 169453 95846 170253 6 dmem_client_request_get[85]
port 95 nsew signal output
rlabel metal2 s 96618 169453 96674 170253 6 dmem_client_request_get[86]
port 96 nsew signal output
rlabel metal2 s 97446 169453 97502 170253 6 dmem_client_request_get[87]
port 97 nsew signal output
rlabel metal2 s 98182 169453 98238 170253 6 dmem_client_request_get[88]
port 98 nsew signal output
rlabel metal2 s 99010 169453 99066 170253 6 dmem_client_request_get[89]
port 99 nsew signal output
rlabel metal2 s 16118 169453 16174 170253 6 dmem_client_request_get[8]
port 100 nsew signal output
rlabel metal2 s 99746 169453 99802 170253 6 dmem_client_request_get[90]
port 101 nsew signal output
rlabel metal2 s 100574 169453 100630 170253 6 dmem_client_request_get[91]
port 102 nsew signal output
rlabel metal2 s 101310 169453 101366 170253 6 dmem_client_request_get[92]
port 103 nsew signal output
rlabel metal2 s 102138 169453 102194 170253 6 dmem_client_request_get[93]
port 104 nsew signal output
rlabel metal2 s 102966 169453 103022 170253 6 dmem_client_request_get[94]
port 105 nsew signal output
rlabel metal2 s 103702 169453 103758 170253 6 dmem_client_request_get[95]
port 106 nsew signal output
rlabel metal2 s 104530 169453 104586 170253 6 dmem_client_request_get[96]
port 107 nsew signal output
rlabel metal2 s 105266 169453 105322 170253 6 dmem_client_request_get[97]
port 108 nsew signal output
rlabel metal2 s 106094 169453 106150 170253 6 dmem_client_request_get[98]
port 109 nsew signal output
rlabel metal2 s 106830 169453 106886 170253 6 dmem_client_request_get[99]
port 110 nsew signal output
rlabel metal2 s 17682 169453 17738 170253 6 dmem_client_request_get[9]
port 111 nsew signal output
rlabel metal2 s 4250 169453 4306 170253 6 dmem_client_response_put[0]
port 112 nsew signal input
rlabel metal2 s 20074 169453 20130 170253 6 dmem_client_response_put[10]
port 113 nsew signal input
rlabel metal2 s 21638 169453 21694 170253 6 dmem_client_response_put[11]
port 114 nsew signal input
rlabel metal2 s 23202 169453 23258 170253 6 dmem_client_response_put[12]
port 115 nsew signal input
rlabel metal2 s 24766 169453 24822 170253 6 dmem_client_response_put[13]
port 116 nsew signal input
rlabel metal2 s 26422 169453 26478 170253 6 dmem_client_response_put[14]
port 117 nsew signal input
rlabel metal2 s 27986 169453 28042 170253 6 dmem_client_response_put[15]
port 118 nsew signal input
rlabel metal2 s 29550 169453 29606 170253 6 dmem_client_response_put[16]
port 119 nsew signal input
rlabel metal2 s 31114 169453 31170 170253 6 dmem_client_response_put[17]
port 120 nsew signal input
rlabel metal2 s 32678 169453 32734 170253 6 dmem_client_response_put[18]
port 121 nsew signal input
rlabel metal2 s 34242 169453 34298 170253 6 dmem_client_response_put[19]
port 122 nsew signal input
rlabel metal2 s 5906 169453 5962 170253 6 dmem_client_response_put[1]
port 123 nsew signal input
rlabel metal2 s 35806 169453 35862 170253 6 dmem_client_response_put[20]
port 124 nsew signal input
rlabel metal2 s 37462 169453 37518 170253 6 dmem_client_response_put[21]
port 125 nsew signal input
rlabel metal2 s 39026 169453 39082 170253 6 dmem_client_response_put[22]
port 126 nsew signal input
rlabel metal2 s 40590 169453 40646 170253 6 dmem_client_response_put[23]
port 127 nsew signal input
rlabel metal2 s 42154 169453 42210 170253 6 dmem_client_response_put[24]
port 128 nsew signal input
rlabel metal2 s 43718 169453 43774 170253 6 dmem_client_response_put[25]
port 129 nsew signal input
rlabel metal2 s 45282 169453 45338 170253 6 dmem_client_response_put[26]
port 130 nsew signal input
rlabel metal2 s 46938 169453 46994 170253 6 dmem_client_response_put[27]
port 131 nsew signal input
rlabel metal2 s 48502 169453 48558 170253 6 dmem_client_response_put[28]
port 132 nsew signal input
rlabel metal2 s 50066 169453 50122 170253 6 dmem_client_response_put[29]
port 133 nsew signal input
rlabel metal2 s 7470 169453 7526 170253 6 dmem_client_response_put[2]
port 134 nsew signal input
rlabel metal2 s 51630 169453 51686 170253 6 dmem_client_response_put[30]
port 135 nsew signal input
rlabel metal2 s 53194 169453 53250 170253 6 dmem_client_response_put[31]
port 136 nsew signal input
rlabel metal2 s 9034 169453 9090 170253 6 dmem_client_response_put[3]
port 137 nsew signal input
rlabel metal2 s 10598 169453 10654 170253 6 dmem_client_response_put[4]
port 138 nsew signal input
rlabel metal2 s 12162 169453 12218 170253 6 dmem_client_response_put[5]
port 139 nsew signal input
rlabel metal2 s 13726 169453 13782 170253 6 dmem_client_response_put[6]
port 140 nsew signal input
rlabel metal2 s 15290 169453 15346 170253 6 dmem_client_response_put[7]
port 141 nsew signal input
rlabel metal2 s 16946 169453 17002 170253 6 dmem_client_response_put[8]
port 142 nsew signal input
rlabel metal2 s 18510 169453 18566 170253 6 dmem_client_response_put[9]
port 143 nsew signal input
rlabel metal2 s 110786 169453 110842 170253 6 imem_client_request_get[0]
port 144 nsew signal output
rlabel metal2 s 126610 169453 126666 170253 6 imem_client_request_get[10]
port 145 nsew signal output
rlabel metal2 s 128174 169453 128230 170253 6 imem_client_request_get[11]
port 146 nsew signal output
rlabel metal2 s 129738 169453 129794 170253 6 imem_client_request_get[12]
port 147 nsew signal output
rlabel metal2 s 131302 169453 131358 170253 6 imem_client_request_get[13]
port 148 nsew signal output
rlabel metal2 s 132958 169453 133014 170253 6 imem_client_request_get[14]
port 149 nsew signal output
rlabel metal2 s 134522 169453 134578 170253 6 imem_client_request_get[15]
port 150 nsew signal output
rlabel metal2 s 136086 169453 136142 170253 6 imem_client_request_get[16]
port 151 nsew signal output
rlabel metal2 s 137650 169453 137706 170253 6 imem_client_request_get[17]
port 152 nsew signal output
rlabel metal2 s 139214 169453 139270 170253 6 imem_client_request_get[18]
port 153 nsew signal output
rlabel metal2 s 140778 169453 140834 170253 6 imem_client_request_get[19]
port 154 nsew signal output
rlabel metal2 s 112442 169453 112498 170253 6 imem_client_request_get[1]
port 155 nsew signal output
rlabel metal2 s 142342 169453 142398 170253 6 imem_client_request_get[20]
port 156 nsew signal output
rlabel metal2 s 143998 169453 144054 170253 6 imem_client_request_get[21]
port 157 nsew signal output
rlabel metal2 s 145562 169453 145618 170253 6 imem_client_request_get[22]
port 158 nsew signal output
rlabel metal2 s 147126 169453 147182 170253 6 imem_client_request_get[23]
port 159 nsew signal output
rlabel metal2 s 148690 169453 148746 170253 6 imem_client_request_get[24]
port 160 nsew signal output
rlabel metal2 s 150254 169453 150310 170253 6 imem_client_request_get[25]
port 161 nsew signal output
rlabel metal2 s 151818 169453 151874 170253 6 imem_client_request_get[26]
port 162 nsew signal output
rlabel metal2 s 153474 169453 153530 170253 6 imem_client_request_get[27]
port 163 nsew signal output
rlabel metal2 s 155038 169453 155094 170253 6 imem_client_request_get[28]
port 164 nsew signal output
rlabel metal2 s 156602 169453 156658 170253 6 imem_client_request_get[29]
port 165 nsew signal output
rlabel metal2 s 114006 169453 114062 170253 6 imem_client_request_get[2]
port 166 nsew signal output
rlabel metal2 s 158166 169453 158222 170253 6 imem_client_request_get[30]
port 167 nsew signal output
rlabel metal2 s 159730 169453 159786 170253 6 imem_client_request_get[31]
port 168 nsew signal output
rlabel metal2 s 115570 169453 115626 170253 6 imem_client_request_get[3]
port 169 nsew signal output
rlabel metal2 s 117134 169453 117190 170253 6 imem_client_request_get[4]
port 170 nsew signal output
rlabel metal2 s 118698 169453 118754 170253 6 imem_client_request_get[5]
port 171 nsew signal output
rlabel metal2 s 120262 169453 120318 170253 6 imem_client_request_get[6]
port 172 nsew signal output
rlabel metal2 s 121826 169453 121882 170253 6 imem_client_request_get[7]
port 173 nsew signal output
rlabel metal2 s 123482 169453 123538 170253 6 imem_client_request_get[8]
port 174 nsew signal output
rlabel metal2 s 125046 169453 125102 170253 6 imem_client_request_get[9]
port 175 nsew signal output
rlabel metal2 s 111614 169453 111670 170253 6 imem_client_response_put[0]
port 176 nsew signal input
rlabel metal2 s 127346 169453 127402 170253 6 imem_client_response_put[10]
port 177 nsew signal input
rlabel metal2 s 129002 169453 129058 170253 6 imem_client_response_put[11]
port 178 nsew signal input
rlabel metal2 s 130566 169453 130622 170253 6 imem_client_response_put[12]
port 179 nsew signal input
rlabel metal2 s 132130 169453 132186 170253 6 imem_client_response_put[13]
port 180 nsew signal input
rlabel metal2 s 133694 169453 133750 170253 6 imem_client_response_put[14]
port 181 nsew signal input
rlabel metal2 s 135258 169453 135314 170253 6 imem_client_response_put[15]
port 182 nsew signal input
rlabel metal2 s 136822 169453 136878 170253 6 imem_client_response_put[16]
port 183 nsew signal input
rlabel metal2 s 138478 169453 138534 170253 6 imem_client_response_put[17]
port 184 nsew signal input
rlabel metal2 s 140042 169453 140098 170253 6 imem_client_response_put[18]
port 185 nsew signal input
rlabel metal2 s 141606 169453 141662 170253 6 imem_client_response_put[19]
port 186 nsew signal input
rlabel metal2 s 113178 169453 113234 170253 6 imem_client_response_put[1]
port 187 nsew signal input
rlabel metal2 s 143170 169453 143226 170253 6 imem_client_response_put[20]
port 188 nsew signal input
rlabel metal2 s 144734 169453 144790 170253 6 imem_client_response_put[21]
port 189 nsew signal input
rlabel metal2 s 146298 169453 146354 170253 6 imem_client_response_put[22]
port 190 nsew signal input
rlabel metal2 s 147862 169453 147918 170253 6 imem_client_response_put[23]
port 191 nsew signal input
rlabel metal2 s 149518 169453 149574 170253 6 imem_client_response_put[24]
port 192 nsew signal input
rlabel metal2 s 151082 169453 151138 170253 6 imem_client_response_put[25]
port 193 nsew signal input
rlabel metal2 s 152646 169453 152702 170253 6 imem_client_response_put[26]
port 194 nsew signal input
rlabel metal2 s 154210 169453 154266 170253 6 imem_client_response_put[27]
port 195 nsew signal input
rlabel metal2 s 155774 169453 155830 170253 6 imem_client_response_put[28]
port 196 nsew signal input
rlabel metal2 s 157338 169453 157394 170253 6 imem_client_response_put[29]
port 197 nsew signal input
rlabel metal2 s 114742 169453 114798 170253 6 imem_client_response_put[2]
port 198 nsew signal input
rlabel metal2 s 158994 169453 159050 170253 6 imem_client_response_put[30]
port 199 nsew signal input
rlabel metal2 s 160558 169453 160614 170253 6 imem_client_response_put[31]
port 200 nsew signal input
rlabel metal2 s 116306 169453 116362 170253 6 imem_client_response_put[3]
port 201 nsew signal input
rlabel metal2 s 117962 169453 118018 170253 6 imem_client_response_put[4]
port 202 nsew signal input
rlabel metal2 s 119526 169453 119582 170253 6 imem_client_response_put[5]
port 203 nsew signal input
rlabel metal2 s 121090 169453 121146 170253 6 imem_client_response_put[6]
port 204 nsew signal input
rlabel metal2 s 122654 169453 122710 170253 6 imem_client_response_put[7]
port 205 nsew signal input
rlabel metal2 s 124218 169453 124274 170253 6 imem_client_response_put[8]
port 206 nsew signal input
rlabel metal2 s 125782 169453 125838 170253 6 imem_client_response_put[9]
port 207 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 readPC[0]
port 208 nsew signal output
rlabel metal3 s 167309 164840 168109 164960 6 readPC[10]
port 209 nsew signal output
rlabel metal2 s 84014 0 84070 800 6 readPC[11]
port 210 nsew signal output
rlabel metal2 s 162858 169453 162914 170253 6 readPC[12]
port 211 nsew signal output
rlabel metal3 s 0 76440 800 76560 6 readPC[13]
port 212 nsew signal output
rlabel metal3 s 167309 166336 168109 166456 6 readPC[14]
port 213 nsew signal output
rlabel metal3 s 0 93576 800 93696 6 readPC[15]
port 214 nsew signal output
rlabel metal2 s 102690 0 102746 800 6 readPC[16]
port 215 nsew signal output
rlabel metal3 s 0 110576 800 110696 6 readPC[17]
port 216 nsew signal output
rlabel metal3 s 167309 167832 168109 167952 6 readPC[18]
port 217 nsew signal output
rlabel metal2 s 163686 169453 163742 170253 6 readPC[19]
port 218 nsew signal output
rlabel metal3 s 0 25440 800 25560 6 readPC[1]
port 219 nsew signal output
rlabel metal2 s 164514 169453 164570 170253 6 readPC[20]
port 220 nsew signal output
rlabel metal2 s 165250 169453 165306 170253 6 readPC[21]
port 221 nsew signal output
rlabel metal3 s 0 127576 800 127696 6 readPC[22]
port 222 nsew signal output
rlabel metal2 s 121366 0 121422 800 6 readPC[23]
port 223 nsew signal output
rlabel metal3 s 0 144576 800 144696 6 readPC[24]
port 224 nsew signal output
rlabel metal2 s 140042 0 140098 800 6 readPC[25]
port 225 nsew signal output
rlabel metal2 s 166078 169453 166134 170253 6 readPC[26]
port 226 nsew signal output
rlabel metal2 s 166814 169453 166870 170253 6 readPC[27]
port 227 nsew signal output
rlabel metal2 s 158718 0 158774 800 6 readPC[28]
port 228 nsew signal output
rlabel metal2 s 167642 169453 167698 170253 6 readPC[29]
port 229 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 readPC[2]
port 230 nsew signal output
rlabel metal3 s 167309 169328 168109 169448 6 readPC[30]
port 231 nsew signal output
rlabel metal3 s 0 161576 800 161696 6 readPC[31]
port 232 nsew signal output
rlabel metal2 s 161294 169453 161350 170253 6 readPC[3]
port 233 nsew signal output
rlabel metal2 s 162122 169453 162178 170253 6 readPC[4]
port 234 nsew signal output
rlabel metal3 s 167309 160352 168109 160472 6 readPC[5]
port 235 nsew signal output
rlabel metal3 s 167309 161848 168109 161968 6 readPC[6]
port 236 nsew signal output
rlabel metal3 s 0 42440 800 42560 6 readPC[7]
port 237 nsew signal output
rlabel metal3 s 0 59440 800 59560 6 readPC[8]
port 238 nsew signal output
rlabel metal3 s 167309 163344 168109 163464 6 readPC[9]
port 239 nsew signal output
rlabel metal3 s 167309 688 168109 808 6 sysmem_client_ack_i
port 240 nsew signal input
rlabel metal3 s 167309 9664 168109 9784 6 sysmem_client_adr_o[0]
port 241 nsew signal output
rlabel metal3 s 167309 60936 168109 61056 6 sysmem_client_adr_o[10]
port 242 nsew signal output
rlabel metal3 s 167309 65424 168109 65544 6 sysmem_client_adr_o[11]
port 243 nsew signal output
rlabel metal3 s 167309 69912 168109 70032 6 sysmem_client_adr_o[12]
port 244 nsew signal output
rlabel metal3 s 167309 74400 168109 74520 6 sysmem_client_adr_o[13]
port 245 nsew signal output
rlabel metal3 s 167309 79024 168109 79144 6 sysmem_client_adr_o[14]
port 246 nsew signal output
rlabel metal3 s 167309 83512 168109 83632 6 sysmem_client_adr_o[15]
port 247 nsew signal output
rlabel metal3 s 167309 88000 168109 88120 6 sysmem_client_adr_o[16]
port 248 nsew signal output
rlabel metal3 s 167309 92488 168109 92608 6 sysmem_client_adr_o[17]
port 249 nsew signal output
rlabel metal3 s 167309 97112 168109 97232 6 sysmem_client_adr_o[18]
port 250 nsew signal output
rlabel metal3 s 167309 101600 168109 101720 6 sysmem_client_adr_o[19]
port 251 nsew signal output
rlabel metal3 s 167309 15648 168109 15768 6 sysmem_client_adr_o[1]
port 252 nsew signal output
rlabel metal3 s 167309 106088 168109 106208 6 sysmem_client_adr_o[20]
port 253 nsew signal output
rlabel metal3 s 167309 110576 168109 110696 6 sysmem_client_adr_o[21]
port 254 nsew signal output
rlabel metal3 s 167309 115200 168109 115320 6 sysmem_client_adr_o[22]
port 255 nsew signal output
rlabel metal3 s 167309 119688 168109 119808 6 sysmem_client_adr_o[23]
port 256 nsew signal output
rlabel metal3 s 167309 124176 168109 124296 6 sysmem_client_adr_o[24]
port 257 nsew signal output
rlabel metal3 s 167309 128664 168109 128784 6 sysmem_client_adr_o[25]
port 258 nsew signal output
rlabel metal3 s 167309 133288 168109 133408 6 sysmem_client_adr_o[26]
port 259 nsew signal output
rlabel metal3 s 167309 137776 168109 137896 6 sysmem_client_adr_o[27]
port 260 nsew signal output
rlabel metal3 s 167309 142264 168109 142384 6 sysmem_client_adr_o[28]
port 261 nsew signal output
rlabel metal3 s 167309 146752 168109 146872 6 sysmem_client_adr_o[29]
port 262 nsew signal output
rlabel metal3 s 167309 21768 168109 21888 6 sysmem_client_adr_o[2]
port 263 nsew signal output
rlabel metal3 s 167309 151240 168109 151360 6 sysmem_client_adr_o[30]
port 264 nsew signal output
rlabel metal3 s 167309 155864 168109 155984 6 sysmem_client_adr_o[31]
port 265 nsew signal output
rlabel metal3 s 167309 27752 168109 27872 6 sysmem_client_adr_o[3]
port 266 nsew signal output
rlabel metal3 s 167309 33736 168109 33856 6 sysmem_client_adr_o[4]
port 267 nsew signal output
rlabel metal3 s 167309 38224 168109 38344 6 sysmem_client_adr_o[5]
port 268 nsew signal output
rlabel metal3 s 167309 42848 168109 42968 6 sysmem_client_adr_o[6]
port 269 nsew signal output
rlabel metal3 s 167309 47336 168109 47456 6 sysmem_client_adr_o[7]
port 270 nsew signal output
rlabel metal3 s 167309 51824 168109 51944 6 sysmem_client_adr_o[8]
port 271 nsew signal output
rlabel metal3 s 167309 56312 168109 56432 6 sysmem_client_adr_o[9]
port 272 nsew signal output
rlabel metal3 s 167309 2184 168109 2304 6 sysmem_client_cyc_o
port 273 nsew signal output
rlabel metal3 s 167309 11160 168109 11280 6 sysmem_client_dat_i[0]
port 274 nsew signal input
rlabel metal3 s 167309 62432 168109 62552 6 sysmem_client_dat_i[10]
port 275 nsew signal input
rlabel metal3 s 167309 66920 168109 67040 6 sysmem_client_dat_i[11]
port 276 nsew signal input
rlabel metal3 s 167309 71408 168109 71528 6 sysmem_client_dat_i[12]
port 277 nsew signal input
rlabel metal3 s 167309 75896 168109 76016 6 sysmem_client_dat_i[13]
port 278 nsew signal input
rlabel metal3 s 167309 80520 168109 80640 6 sysmem_client_dat_i[14]
port 279 nsew signal input
rlabel metal3 s 167309 85008 168109 85128 6 sysmem_client_dat_i[15]
port 280 nsew signal input
rlabel metal3 s 167309 89496 168109 89616 6 sysmem_client_dat_i[16]
port 281 nsew signal input
rlabel metal3 s 167309 93984 168109 94104 6 sysmem_client_dat_i[17]
port 282 nsew signal input
rlabel metal3 s 167309 98608 168109 98728 6 sysmem_client_dat_i[18]
port 283 nsew signal input
rlabel metal3 s 167309 103096 168109 103216 6 sysmem_client_dat_i[19]
port 284 nsew signal input
rlabel metal3 s 167309 17144 168109 17264 6 sysmem_client_dat_i[1]
port 285 nsew signal input
rlabel metal3 s 167309 107584 168109 107704 6 sysmem_client_dat_i[20]
port 286 nsew signal input
rlabel metal3 s 167309 112072 168109 112192 6 sysmem_client_dat_i[21]
port 287 nsew signal input
rlabel metal3 s 167309 116696 168109 116816 6 sysmem_client_dat_i[22]
port 288 nsew signal input
rlabel metal3 s 167309 121184 168109 121304 6 sysmem_client_dat_i[23]
port 289 nsew signal input
rlabel metal3 s 167309 125672 168109 125792 6 sysmem_client_dat_i[24]
port 290 nsew signal input
rlabel metal3 s 167309 130160 168109 130280 6 sysmem_client_dat_i[25]
port 291 nsew signal input
rlabel metal3 s 167309 134784 168109 134904 6 sysmem_client_dat_i[26]
port 292 nsew signal input
rlabel metal3 s 167309 139272 168109 139392 6 sysmem_client_dat_i[27]
port 293 nsew signal input
rlabel metal3 s 167309 143760 168109 143880 6 sysmem_client_dat_i[28]
port 294 nsew signal input
rlabel metal3 s 167309 148248 168109 148368 6 sysmem_client_dat_i[29]
port 295 nsew signal input
rlabel metal3 s 167309 23264 168109 23384 6 sysmem_client_dat_i[2]
port 296 nsew signal input
rlabel metal3 s 167309 152872 168109 152992 6 sysmem_client_dat_i[30]
port 297 nsew signal input
rlabel metal3 s 167309 157360 168109 157480 6 sysmem_client_dat_i[31]
port 298 nsew signal input
rlabel metal3 s 167309 29248 168109 29368 6 sysmem_client_dat_i[3]
port 299 nsew signal input
rlabel metal3 s 167309 35232 168109 35352 6 sysmem_client_dat_i[4]
port 300 nsew signal input
rlabel metal3 s 167309 39856 168109 39976 6 sysmem_client_dat_i[5]
port 301 nsew signal input
rlabel metal3 s 167309 44344 168109 44464 6 sysmem_client_dat_i[6]
port 302 nsew signal input
rlabel metal3 s 167309 48832 168109 48952 6 sysmem_client_dat_i[7]
port 303 nsew signal input
rlabel metal3 s 167309 53320 168109 53440 6 sysmem_client_dat_i[8]
port 304 nsew signal input
rlabel metal3 s 167309 57944 168109 58064 6 sysmem_client_dat_i[9]
port 305 nsew signal input
rlabel metal3 s 167309 12656 168109 12776 6 sysmem_client_dat_o[0]
port 306 nsew signal output
rlabel metal3 s 167309 63928 168109 64048 6 sysmem_client_dat_o[10]
port 307 nsew signal output
rlabel metal3 s 167309 68416 168109 68536 6 sysmem_client_dat_o[11]
port 308 nsew signal output
rlabel metal3 s 167309 72904 168109 73024 6 sysmem_client_dat_o[12]
port 309 nsew signal output
rlabel metal3 s 167309 77528 168109 77648 6 sysmem_client_dat_o[13]
port 310 nsew signal output
rlabel metal3 s 167309 82016 168109 82136 6 sysmem_client_dat_o[14]
port 311 nsew signal output
rlabel metal3 s 167309 86504 168109 86624 6 sysmem_client_dat_o[15]
port 312 nsew signal output
rlabel metal3 s 167309 90992 168109 91112 6 sysmem_client_dat_o[16]
port 313 nsew signal output
rlabel metal3 s 167309 95616 168109 95736 6 sysmem_client_dat_o[17]
port 314 nsew signal output
rlabel metal3 s 167309 100104 168109 100224 6 sysmem_client_dat_o[18]
port 315 nsew signal output
rlabel metal3 s 167309 104592 168109 104712 6 sysmem_client_dat_o[19]
port 316 nsew signal output
rlabel metal3 s 167309 18640 168109 18760 6 sysmem_client_dat_o[1]
port 317 nsew signal output
rlabel metal3 s 167309 109080 168109 109200 6 sysmem_client_dat_o[20]
port 318 nsew signal output
rlabel metal3 s 167309 113568 168109 113688 6 sysmem_client_dat_o[21]
port 319 nsew signal output
rlabel metal3 s 167309 118192 168109 118312 6 sysmem_client_dat_o[22]
port 320 nsew signal output
rlabel metal3 s 167309 122680 168109 122800 6 sysmem_client_dat_o[23]
port 321 nsew signal output
rlabel metal3 s 167309 127168 168109 127288 6 sysmem_client_dat_o[24]
port 322 nsew signal output
rlabel metal3 s 167309 131656 168109 131776 6 sysmem_client_dat_o[25]
port 323 nsew signal output
rlabel metal3 s 167309 136280 168109 136400 6 sysmem_client_dat_o[26]
port 324 nsew signal output
rlabel metal3 s 167309 140768 168109 140888 6 sysmem_client_dat_o[27]
port 325 nsew signal output
rlabel metal3 s 167309 145256 168109 145376 6 sysmem_client_dat_o[28]
port 326 nsew signal output
rlabel metal3 s 167309 149744 168109 149864 6 sysmem_client_dat_o[29]
port 327 nsew signal output
rlabel metal3 s 167309 24760 168109 24880 6 sysmem_client_dat_o[2]
port 328 nsew signal output
rlabel metal3 s 167309 154368 168109 154488 6 sysmem_client_dat_o[30]
port 329 nsew signal output
rlabel metal3 s 167309 158856 168109 158976 6 sysmem_client_dat_o[31]
port 330 nsew signal output
rlabel metal3 s 167309 30744 168109 30864 6 sysmem_client_dat_o[3]
port 331 nsew signal output
rlabel metal3 s 167309 36728 168109 36848 6 sysmem_client_dat_o[4]
port 332 nsew signal output
rlabel metal3 s 167309 41352 168109 41472 6 sysmem_client_dat_o[5]
port 333 nsew signal output
rlabel metal3 s 167309 45840 168109 45960 6 sysmem_client_dat_o[6]
port 334 nsew signal output
rlabel metal3 s 167309 50328 168109 50448 6 sysmem_client_dat_o[7]
port 335 nsew signal output
rlabel metal3 s 167309 54816 168109 54936 6 sysmem_client_dat_o[8]
port 336 nsew signal output
rlabel metal3 s 167309 59440 168109 59560 6 sysmem_client_dat_o[9]
port 337 nsew signal output
rlabel metal3 s 167309 3680 168109 3800 6 sysmem_client_err_i
port 338 nsew signal input
rlabel metal3 s 167309 5176 168109 5296 6 sysmem_client_rty_i
port 339 nsew signal input
rlabel metal3 s 167309 14152 168109 14272 6 sysmem_client_sel_o[0]
port 340 nsew signal output
rlabel metal3 s 167309 20272 168109 20392 6 sysmem_client_sel_o[1]
port 341 nsew signal output
rlabel metal3 s 167309 26256 168109 26376 6 sysmem_client_sel_o[2]
port 342 nsew signal output
rlabel metal3 s 167309 32240 168109 32360 6 sysmem_client_sel_o[3]
port 343 nsew signal output
rlabel metal3 s 167309 6672 168109 6792 6 sysmem_client_stb_o
port 344 nsew signal output
rlabel metal3 s 167309 8168 168109 8288 6 sysmem_client_we_o
port 345 nsew signal output
rlabel metal4 s 4208 2128 4528 167600 6 vccd1
port 346 nsew power input
rlabel metal4 s 34928 2128 35248 167600 6 vccd1
port 346 nsew power input
rlabel metal4 s 65648 2128 65968 167600 6 vccd1
port 346 nsew power input
rlabel metal4 s 96368 2128 96688 167600 6 vccd1
port 346 nsew power input
rlabel metal4 s 127088 2128 127408 167600 6 vccd1
port 346 nsew power input
rlabel metal4 s 157808 2128 158128 167600 6 vccd1
port 346 nsew power input
rlabel metal4 s 19568 2128 19888 167600 6 vssd1
port 347 nsew ground input
rlabel metal4 s 50288 2128 50608 167600 6 vssd1
port 347 nsew ground input
rlabel metal4 s 81008 2128 81328 167600 6 vssd1
port 347 nsew ground input
rlabel metal4 s 111728 2128 112048 167600 6 vssd1
port 347 nsew ground input
rlabel metal4 s 142448 2128 142768 167600 6 vssd1
port 347 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 168109 170253
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 73598818
string GDS_FILE /home/q3k/sky130/qf105/openlane/mkLanaiCPU/runs/mkLanaiCPU/results/finishing/mkLanaiCPU.magic.gds
string GDS_START 1597022
<< end >>

