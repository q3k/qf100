VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mkLanaiCPU
  CLASS BLOCK ;
  FOREIGN mkLanaiCPU ;
  ORIGIN 0.000 0.000 ;
  SIZE 839.870 BY 850.590 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 773.880 839.870 774.480 ;
    END
  END CLK
  PIN EN_dmem_client_request_get
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 846.590 2.210 850.590 ;
    END
  END EN_dmem_client_request_get
  PIN EN_dmem_client_response_put
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 846.590 5.890 850.590 ;
    END
  END EN_dmem_client_response_put
  PIN EN_imem_client_request_get
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 846.590 545.930 850.590 ;
    END
  END EN_imem_client_request_get
  PIN EN_imem_client_response_put
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 846.590 550.070 850.590 ;
    END
  END EN_imem_client_response_put
  PIN RDY_dmem_client_request_get
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 846.590 10.030 850.590 ;
    END
  END RDY_dmem_client_request_get
  PIN RDY_dmem_client_response_put
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 846.590 14.170 850.590 ;
    END
  END RDY_dmem_client_response_put
  PIN RDY_imem_client_request_get
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 846.590 553.750 850.590 ;
    END
  END RDY_imem_client_request_get
  PIN RDY_imem_client_response_put
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 846.590 557.890 850.590 ;
    END
  END RDY_imem_client_response_put
  PIN RDY_readPC
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END RDY_readPC
  PIN RST_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END RST_N
  PIN dmem_client_request_get[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 846.590 17.850 850.590 ;
    END
  END dmem_client_request_get[0]
  PIN dmem_client_request_get[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 846.590 97.890 850.590 ;
    END
  END dmem_client_request_get[10]
  PIN dmem_client_request_get[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 846.590 106.170 850.590 ;
    END
  END dmem_client_request_get[11]
  PIN dmem_client_request_get[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 846.590 113.990 850.590 ;
    END
  END dmem_client_request_get[12]
  PIN dmem_client_request_get[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 846.590 121.810 850.590 ;
    END
  END dmem_client_request_get[13]
  PIN dmem_client_request_get[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 846.590 130.090 850.590 ;
    END
  END dmem_client_request_get[14]
  PIN dmem_client_request_get[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 846.590 137.910 850.590 ;
    END
  END dmem_client_request_get[15]
  PIN dmem_client_request_get[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 846.590 146.190 850.590 ;
    END
  END dmem_client_request_get[16]
  PIN dmem_client_request_get[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 846.590 154.010 850.590 ;
    END
  END dmem_client_request_get[17]
  PIN dmem_client_request_get[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 846.590 161.830 850.590 ;
    END
  END dmem_client_request_get[18]
  PIN dmem_client_request_get[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 846.590 170.110 850.590 ;
    END
  END dmem_client_request_get[19]
  PIN dmem_client_request_get[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 846.590 26.130 850.590 ;
    END
  END dmem_client_request_get[1]
  PIN dmem_client_request_get[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 846.590 177.930 850.590 ;
    END
  END dmem_client_request_get[20]
  PIN dmem_client_request_get[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 846.590 185.750 850.590 ;
    END
  END dmem_client_request_get[21]
  PIN dmem_client_request_get[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 846.590 194.030 850.590 ;
    END
  END dmem_client_request_get[22]
  PIN dmem_client_request_get[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 846.590 201.850 850.590 ;
    END
  END dmem_client_request_get[23]
  PIN dmem_client_request_get[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 846.590 210.130 850.590 ;
    END
  END dmem_client_request_get[24]
  PIN dmem_client_request_get[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 846.590 217.950 850.590 ;
    END
  END dmem_client_request_get[25]
  PIN dmem_client_request_get[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 846.590 225.770 850.590 ;
    END
  END dmem_client_request_get[26]
  PIN dmem_client_request_get[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 846.590 234.050 850.590 ;
    END
  END dmem_client_request_get[27]
  PIN dmem_client_request_get[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 846.590 241.870 850.590 ;
    END
  END dmem_client_request_get[28]
  PIN dmem_client_request_get[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 846.590 250.150 850.590 ;
    END
  END dmem_client_request_get[29]
  PIN dmem_client_request_get[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 846.590 33.950 850.590 ;
    END
  END dmem_client_request_get[2]
  PIN dmem_client_request_get[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 846.590 257.970 850.590 ;
    END
  END dmem_client_request_get[30]
  PIN dmem_client_request_get[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 846.590 265.790 850.590 ;
    END
  END dmem_client_request_get[31]
  PIN dmem_client_request_get[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 846.590 274.070 850.590 ;
    END
  END dmem_client_request_get[32]
  PIN dmem_client_request_get[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 846.590 277.750 850.590 ;
    END
  END dmem_client_request_get[33]
  PIN dmem_client_request_get[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 846.590 281.890 850.590 ;
    END
  END dmem_client_request_get[34]
  PIN dmem_client_request_get[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 846.590 286.030 850.590 ;
    END
  END dmem_client_request_get[35]
  PIN dmem_client_request_get[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 846.590 290.170 850.590 ;
    END
  END dmem_client_request_get[36]
  PIN dmem_client_request_get[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 846.590 293.850 850.590 ;
    END
  END dmem_client_request_get[37]
  PIN dmem_client_request_get[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 846.590 297.990 850.590 ;
    END
  END dmem_client_request_get[38]
  PIN dmem_client_request_get[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 846.590 302.130 850.590 ;
    END
  END dmem_client_request_get[39]
  PIN dmem_client_request_get[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 846.590 41.770 850.590 ;
    END
  END dmem_client_request_get[3]
  PIN dmem_client_request_get[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 846.590 305.810 850.590 ;
    END
  END dmem_client_request_get[40]
  PIN dmem_client_request_get[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 846.590 309.950 850.590 ;
    END
  END dmem_client_request_get[41]
  PIN dmem_client_request_get[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 846.590 314.090 850.590 ;
    END
  END dmem_client_request_get[42]
  PIN dmem_client_request_get[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 846.590 317.770 850.590 ;
    END
  END dmem_client_request_get[43]
  PIN dmem_client_request_get[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 846.590 321.910 850.590 ;
    END
  END dmem_client_request_get[44]
  PIN dmem_client_request_get[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 846.590 326.050 850.590 ;
    END
  END dmem_client_request_get[45]
  PIN dmem_client_request_get[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 846.590 330.190 850.590 ;
    END
  END dmem_client_request_get[46]
  PIN dmem_client_request_get[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 846.590 333.870 850.590 ;
    END
  END dmem_client_request_get[47]
  PIN dmem_client_request_get[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 846.590 338.010 850.590 ;
    END
  END dmem_client_request_get[48]
  PIN dmem_client_request_get[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 846.590 342.150 850.590 ;
    END
  END dmem_client_request_get[49]
  PIN dmem_client_request_get[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 846.590 50.050 850.590 ;
    END
  END dmem_client_request_get[4]
  PIN dmem_client_request_get[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 846.590 345.830 850.590 ;
    END
  END dmem_client_request_get[50]
  PIN dmem_client_request_get[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 846.590 349.970 850.590 ;
    END
  END dmem_client_request_get[51]
  PIN dmem_client_request_get[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 846.590 354.110 850.590 ;
    END
  END dmem_client_request_get[52]
  PIN dmem_client_request_get[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 846.590 357.790 850.590 ;
    END
  END dmem_client_request_get[53]
  PIN dmem_client_request_get[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 846.590 361.930 850.590 ;
    END
  END dmem_client_request_get[54]
  PIN dmem_client_request_get[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 846.590 366.070 850.590 ;
    END
  END dmem_client_request_get[55]
  PIN dmem_client_request_get[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 846.590 369.750 850.590 ;
    END
  END dmem_client_request_get[56]
  PIN dmem_client_request_get[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 846.590 373.890 850.590 ;
    END
  END dmem_client_request_get[57]
  PIN dmem_client_request_get[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 846.590 378.030 850.590 ;
    END
  END dmem_client_request_get[58]
  PIN dmem_client_request_get[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 846.590 382.170 850.590 ;
    END
  END dmem_client_request_get[59]
  PIN dmem_client_request_get[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 846.590 57.870 850.590 ;
    END
  END dmem_client_request_get[5]
  PIN dmem_client_request_get[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 846.590 385.850 850.590 ;
    END
  END dmem_client_request_get[60]
  PIN dmem_client_request_get[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 846.590 389.990 850.590 ;
    END
  END dmem_client_request_get[61]
  PIN dmem_client_request_get[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 846.590 394.130 850.590 ;
    END
  END dmem_client_request_get[62]
  PIN dmem_client_request_get[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 846.590 397.810 850.590 ;
    END
  END dmem_client_request_get[63]
  PIN dmem_client_request_get[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 846.590 401.950 850.590 ;
    END
  END dmem_client_request_get[64]
  PIN dmem_client_request_get[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 846.590 406.090 850.590 ;
    END
  END dmem_client_request_get[65]
  PIN dmem_client_request_get[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 846.590 409.770 850.590 ;
    END
  END dmem_client_request_get[66]
  PIN dmem_client_request_get[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 846.590 413.910 850.590 ;
    END
  END dmem_client_request_get[67]
  PIN dmem_client_request_get[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 846.590 418.050 850.590 ;
    END
  END dmem_client_request_get[68]
  PIN dmem_client_request_get[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 846.590 422.190 850.590 ;
    END
  END dmem_client_request_get[69]
  PIN dmem_client_request_get[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 846.590 66.150 850.590 ;
    END
  END dmem_client_request_get[6]
  PIN dmem_client_request_get[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 846.590 425.870 850.590 ;
    END
  END dmem_client_request_get[70]
  PIN dmem_client_request_get[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 846.590 430.010 850.590 ;
    END
  END dmem_client_request_get[71]
  PIN dmem_client_request_get[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 846.590 434.150 850.590 ;
    END
  END dmem_client_request_get[72]
  PIN dmem_client_request_get[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 846.590 437.830 850.590 ;
    END
  END dmem_client_request_get[73]
  PIN dmem_client_request_get[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 846.590 441.970 850.590 ;
    END
  END dmem_client_request_get[74]
  PIN dmem_client_request_get[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 846.590 446.110 850.590 ;
    END
  END dmem_client_request_get[75]
  PIN dmem_client_request_get[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 846.590 449.790 850.590 ;
    END
  END dmem_client_request_get[76]
  PIN dmem_client_request_get[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 846.590 453.930 850.590 ;
    END
  END dmem_client_request_get[77]
  PIN dmem_client_request_get[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 846.590 458.070 850.590 ;
    END
  END dmem_client_request_get[78]
  PIN dmem_client_request_get[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 846.590 461.750 850.590 ;
    END
  END dmem_client_request_get[79]
  PIN dmem_client_request_get[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 846.590 73.970 850.590 ;
    END
  END dmem_client_request_get[7]
  PIN dmem_client_request_get[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 846.590 465.890 850.590 ;
    END
  END dmem_client_request_get[80]
  PIN dmem_client_request_get[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 846.590 470.030 850.590 ;
    END
  END dmem_client_request_get[81]
  PIN dmem_client_request_get[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 846.590 474.170 850.590 ;
    END
  END dmem_client_request_get[82]
  PIN dmem_client_request_get[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.570 846.590 477.850 850.590 ;
    END
  END dmem_client_request_get[83]
  PIN dmem_client_request_get[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 846.590 481.990 850.590 ;
    END
  END dmem_client_request_get[84]
  PIN dmem_client_request_get[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 846.590 486.130 850.590 ;
    END
  END dmem_client_request_get[85]
  PIN dmem_client_request_get[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 846.590 489.810 850.590 ;
    END
  END dmem_client_request_get[86]
  PIN dmem_client_request_get[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.670 846.590 493.950 850.590 ;
    END
  END dmem_client_request_get[87]
  PIN dmem_client_request_get[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.810 846.590 498.090 850.590 ;
    END
  END dmem_client_request_get[88]
  PIN dmem_client_request_get[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.490 846.590 501.770 850.590 ;
    END
  END dmem_client_request_get[89]
  PIN dmem_client_request_get[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 846.590 81.790 850.590 ;
    END
  END dmem_client_request_get[8]
  PIN dmem_client_request_get[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 846.590 505.910 850.590 ;
    END
  END dmem_client_request_get[90]
  PIN dmem_client_request_get[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 846.590 510.050 850.590 ;
    END
  END dmem_client_request_get[91]
  PIN dmem_client_request_get[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 846.590 513.730 850.590 ;
    END
  END dmem_client_request_get[92]
  PIN dmem_client_request_get[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 846.590 517.870 850.590 ;
    END
  END dmem_client_request_get[93]
  PIN dmem_client_request_get[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 846.590 522.010 850.590 ;
    END
  END dmem_client_request_get[94]
  PIN dmem_client_request_get[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.870 846.590 526.150 850.590 ;
    END
  END dmem_client_request_get[95]
  PIN dmem_client_request_get[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 846.590 529.830 850.590 ;
    END
  END dmem_client_request_get[96]
  PIN dmem_client_request_get[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 846.590 533.970 850.590 ;
    END
  END dmem_client_request_get[97]
  PIN dmem_client_request_get[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 846.590 538.110 850.590 ;
    END
  END dmem_client_request_get[98]
  PIN dmem_client_request_get[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 846.590 541.790 850.590 ;
    END
  END dmem_client_request_get[99]
  PIN dmem_client_request_get[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 846.590 90.070 850.590 ;
    END
  END dmem_client_request_get[9]
  PIN dmem_client_response_put[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 846.590 21.990 850.590 ;
    END
  END dmem_client_response_put[0]
  PIN dmem_client_response_put[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 846.590 102.030 850.590 ;
    END
  END dmem_client_response_put[10]
  PIN dmem_client_response_put[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 846.590 109.850 850.590 ;
    END
  END dmem_client_response_put[11]
  PIN dmem_client_response_put[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 846.590 118.130 850.590 ;
    END
  END dmem_client_response_put[12]
  PIN dmem_client_response_put[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 846.590 125.950 850.590 ;
    END
  END dmem_client_response_put[13]
  PIN dmem_client_response_put[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 846.590 133.770 850.590 ;
    END
  END dmem_client_response_put[14]
  PIN dmem_client_response_put[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 846.590 142.050 850.590 ;
    END
  END dmem_client_response_put[15]
  PIN dmem_client_response_put[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 846.590 149.870 850.590 ;
    END
  END dmem_client_response_put[16]
  PIN dmem_client_response_put[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 846.590 158.150 850.590 ;
    END
  END dmem_client_response_put[17]
  PIN dmem_client_response_put[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 846.590 165.970 850.590 ;
    END
  END dmem_client_response_put[18]
  PIN dmem_client_response_put[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 846.590 173.790 850.590 ;
    END
  END dmem_client_response_put[19]
  PIN dmem_client_response_put[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 846.590 29.810 850.590 ;
    END
  END dmem_client_response_put[1]
  PIN dmem_client_response_put[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 846.590 182.070 850.590 ;
    END
  END dmem_client_response_put[20]
  PIN dmem_client_response_put[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 846.590 189.890 850.590 ;
    END
  END dmem_client_response_put[21]
  PIN dmem_client_response_put[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 846.590 198.170 850.590 ;
    END
  END dmem_client_response_put[22]
  PIN dmem_client_response_put[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 846.590 205.990 850.590 ;
    END
  END dmem_client_response_put[23]
  PIN dmem_client_response_put[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 846.590 213.810 850.590 ;
    END
  END dmem_client_response_put[24]
  PIN dmem_client_response_put[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 846.590 222.090 850.590 ;
    END
  END dmem_client_response_put[25]
  PIN dmem_client_response_put[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 846.590 229.910 850.590 ;
    END
  END dmem_client_response_put[26]
  PIN dmem_client_response_put[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 846.590 238.190 850.590 ;
    END
  END dmem_client_response_put[27]
  PIN dmem_client_response_put[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 846.590 246.010 850.590 ;
    END
  END dmem_client_response_put[28]
  PIN dmem_client_response_put[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 846.590 253.830 850.590 ;
    END
  END dmem_client_response_put[29]
  PIN dmem_client_response_put[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 846.590 38.090 850.590 ;
    END
  END dmem_client_response_put[2]
  PIN dmem_client_response_put[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 846.590 262.110 850.590 ;
    END
  END dmem_client_response_put[30]
  PIN dmem_client_response_put[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 846.590 269.930 850.590 ;
    END
  END dmem_client_response_put[31]
  PIN dmem_client_response_put[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 846.590 45.910 850.590 ;
    END
  END dmem_client_response_put[3]
  PIN dmem_client_response_put[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 846.590 54.190 850.590 ;
    END
  END dmem_client_response_put[4]
  PIN dmem_client_response_put[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 846.590 62.010 850.590 ;
    END
  END dmem_client_response_put[5]
  PIN dmem_client_response_put[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 846.590 69.830 850.590 ;
    END
  END dmem_client_response_put[6]
  PIN dmem_client_response_put[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 846.590 78.110 850.590 ;
    END
  END dmem_client_response_put[7]
  PIN dmem_client_response_put[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 846.590 85.930 850.590 ;
    END
  END dmem_client_response_put[8]
  PIN dmem_client_response_put[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 846.590 93.750 850.590 ;
    END
  END dmem_client_response_put[9]
  PIN imem_client_request_get[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 846.590 562.030 850.590 ;
    END
  END imem_client_request_get[0]
  PIN imem_client_request_get[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 846.590 642.070 850.590 ;
    END
  END imem_client_request_get[10]
  PIN imem_client_request_get[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 846.590 649.890 850.590 ;
    END
  END imem_client_request_get[11]
  PIN imem_client_request_get[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 846.590 658.170 850.590 ;
    END
  END imem_client_request_get[12]
  PIN imem_client_request_get[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.710 846.590 665.990 850.590 ;
    END
  END imem_client_request_get[13]
  PIN imem_client_request_get[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 846.590 673.810 850.590 ;
    END
  END imem_client_request_get[14]
  PIN imem_client_request_get[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 846.590 682.090 850.590 ;
    END
  END imem_client_request_get[15]
  PIN imem_client_request_get[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.630 846.590 689.910 850.590 ;
    END
  END imem_client_request_get[16]
  PIN imem_client_request_get[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 846.590 697.730 850.590 ;
    END
  END imem_client_request_get[17]
  PIN imem_client_request_get[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.730 846.590 706.010 850.590 ;
    END
  END imem_client_request_get[18]
  PIN imem_client_request_get[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.550 846.590 713.830 850.590 ;
    END
  END imem_client_request_get[19]
  PIN imem_client_request_get[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 846.590 569.850 850.590 ;
    END
  END imem_client_request_get[1]
  PIN imem_client_request_get[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.830 846.590 722.110 850.590 ;
    END
  END imem_client_request_get[20]
  PIN imem_client_request_get[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 846.590 729.930 850.590 ;
    END
  END imem_client_request_get[21]
  PIN imem_client_request_get[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 846.590 737.750 850.590 ;
    END
  END imem_client_request_get[22]
  PIN imem_client_request_get[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.750 846.590 746.030 850.590 ;
    END
  END imem_client_request_get[23]
  PIN imem_client_request_get[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 846.590 753.850 850.590 ;
    END
  END imem_client_request_get[24]
  PIN imem_client_request_get[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.850 846.590 762.130 850.590 ;
    END
  END imem_client_request_get[25]
  PIN imem_client_request_get[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 846.590 769.950 850.590 ;
    END
  END imem_client_request_get[26]
  PIN imem_client_request_get[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.490 846.590 777.770 850.590 ;
    END
  END imem_client_request_get[27]
  PIN imem_client_request_get[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 846.590 786.050 850.590 ;
    END
  END imem_client_request_get[28]
  PIN imem_client_request_get[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 846.590 793.870 850.590 ;
    END
  END imem_client_request_get[29]
  PIN imem_client_request_get[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 846.590 578.130 850.590 ;
    END
  END imem_client_request_get[2]
  PIN imem_client_request_get[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 846.590 802.150 850.590 ;
    END
  END imem_client_request_get[30]
  PIN imem_client_request_get[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 846.590 809.970 850.590 ;
    END
  END imem_client_request_get[31]
  PIN imem_client_request_get[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 846.590 585.950 850.590 ;
    END
  END imem_client_request_get[3]
  PIN imem_client_request_get[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 846.590 593.770 850.590 ;
    END
  END imem_client_request_get[4]
  PIN imem_client_request_get[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.770 846.590 602.050 850.590 ;
    END
  END imem_client_request_get[5]
  PIN imem_client_request_get[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 846.590 609.870 850.590 ;
    END
  END imem_client_request_get[6]
  PIN imem_client_request_get[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 846.590 618.150 850.590 ;
    END
  END imem_client_request_get[7]
  PIN imem_client_request_get[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 846.590 625.970 850.590 ;
    END
  END imem_client_request_get[8]
  PIN imem_client_request_get[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.510 846.590 633.790 850.590 ;
    END
  END imem_client_request_get[9]
  PIN imem_client_response_put[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 846.590 566.170 850.590 ;
    END
  END imem_client_response_put[0]
  PIN imem_client_response_put[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.470 846.590 645.750 850.590 ;
    END
  END imem_client_response_put[10]
  PIN imem_client_response_put[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 846.590 654.030 850.590 ;
    END
  END imem_client_response_put[11]
  PIN imem_client_response_put[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.570 846.590 661.850 850.590 ;
    END
  END imem_client_response_put[12]
  PIN imem_client_response_put[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 846.590 670.130 850.590 ;
    END
  END imem_client_response_put[13]
  PIN imem_client_response_put[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.670 846.590 677.950 850.590 ;
    END
  END imem_client_response_put[14]
  PIN imem_client_response_put[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 846.590 685.770 850.590 ;
    END
  END imem_client_response_put[15]
  PIN imem_client_response_put[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 846.590 694.050 850.590 ;
    END
  END imem_client_response_put[16]
  PIN imem_client_response_put[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.590 846.590 701.870 850.590 ;
    END
  END imem_client_response_put[17]
  PIN imem_client_response_put[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.870 846.590 710.150 850.590 ;
    END
  END imem_client_response_put[18]
  PIN imem_client_response_put[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 846.590 717.970 850.590 ;
    END
  END imem_client_response_put[19]
  PIN imem_client_response_put[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 846.590 573.990 850.590 ;
    END
  END imem_client_response_put[1]
  PIN imem_client_response_put[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.510 846.590 725.790 850.590 ;
    END
  END imem_client_response_put[20]
  PIN imem_client_response_put[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.790 846.590 734.070 850.590 ;
    END
  END imem_client_response_put[21]
  PIN imem_client_response_put[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 846.590 741.890 850.590 ;
    END
  END imem_client_response_put[22]
  PIN imem_client_response_put[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 846.590 750.170 850.590 ;
    END
  END imem_client_response_put[23]
  PIN imem_client_response_put[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.710 846.590 757.990 850.590 ;
    END
  END imem_client_response_put[24]
  PIN imem_client_response_put[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 846.590 765.810 850.590 ;
    END
  END imem_client_response_put[25]
  PIN imem_client_response_put[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.810 846.590 774.090 850.590 ;
    END
  END imem_client_response_put[26]
  PIN imem_client_response_put[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.630 846.590 781.910 850.590 ;
    END
  END imem_client_response_put[27]
  PIN imem_client_response_put[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 846.590 789.730 850.590 ;
    END
  END imem_client_response_put[28]
  PIN imem_client_response_put[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 846.590 798.010 850.590 ;
    END
  END imem_client_response_put[29]
  PIN imem_client_response_put[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 846.590 581.810 850.590 ;
    END
  END imem_client_response_put[2]
  PIN imem_client_response_put[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 846.590 805.830 850.590 ;
    END
  END imem_client_response_put[30]
  PIN imem_client_response_put[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.830 846.590 814.110 850.590 ;
    END
  END imem_client_response_put[31]
  PIN imem_client_response_put[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 846.590 590.090 850.590 ;
    END
  END imem_client_response_put[3]
  PIN imem_client_response_put[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 846.590 597.910 850.590 ;
    END
  END imem_client_response_put[4]
  PIN imem_client_response_put[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 846.590 605.730 850.590 ;
    END
  END imem_client_response_put[5]
  PIN imem_client_response_put[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.730 846.590 614.010 850.590 ;
    END
  END imem_client_response_put[6]
  PIN imem_client_response_put[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 846.590 621.830 850.590 ;
    END
  END imem_client_response_put[7]
  PIN imem_client_response_put[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 846.590 630.110 850.590 ;
    END
  END imem_client_response_put[8]
  PIN imem_client_response_put[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 846.590 637.930 850.590 ;
    END
  END imem_client_response_put[9]
  PIN readPC[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 781.360 839.870 781.960 ;
    END
  END readPC[0]
  PIN readPC[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END readPC[10]
  PIN readPC[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.790 846.590 826.070 850.590 ;
    END
  END readPC[11]
  PIN readPC[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 809.920 839.870 810.520 ;
    END
  END readPC[12]
  PIN readPC[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.470 846.590 829.750 850.590 ;
    END
  END readPC[13]
  PIN readPC[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 4.000 294.400 ;
    END
  END readPC[14]
  PIN readPC[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.610 846.590 833.890 850.590 ;
    END
  END readPC[15]
  PIN readPC[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 817.400 839.870 818.000 ;
    END
  END readPC[16]
  PIN readPC[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 824.880 839.870 825.480 ;
    END
  END readPC[17]
  PIN readPC[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.760 4.000 360.360 ;
    END
  END readPC[18]
  PIN readPC[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END readPC[19]
  PIN readPC[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 788.160 839.870 788.760 ;
    END
  END readPC[1]
  PIN readPC[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 0.000 587.790 4.000 ;
    END
  END readPC[20]
  PIN readPC[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 490.320 4.000 490.920 ;
    END
  END readPC[21]
  PIN readPC[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 831.680 839.870 832.280 ;
    END
  END readPC[22]
  PIN readPC[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.410 0.000 755.690 4.000 ;
    END
  END readPC[23]
  PIN readPC[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 839.160 839.870 839.760 ;
    END
  END readPC[24]
  PIN readPC[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 555.600 4.000 556.200 ;
    END
  END readPC[25]
  PIN readPC[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 621.560 4.000 622.160 ;
    END
  END readPC[26]
  PIN readPC[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END readPC[27]
  PIN readPC[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 846.640 839.870 847.240 ;
    END
  END readPC[28]
  PIN readPC[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.750 846.590 838.030 850.590 ;
    END
  END readPC[29]
  PIN readPC[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 795.640 839.870 796.240 ;
    END
  END readPC[2]
  PIN readPC[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.120 4.000 752.720 ;
    END
  END readPC[30]
  PIN readPC[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 817.400 4.000 818.000 ;
    END
  END readPC[31]
  PIN readPC[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 803.120 839.870 803.720 ;
    END
  END readPC[3]
  PIN readPC[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END readPC[4]
  PIN readPC[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END readPC[5]
  PIN readPC[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END readPC[6]
  PIN readPC[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END readPC[7]
  PIN readPC[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.510 846.590 817.790 850.590 ;
    END
  END readPC[8]
  PIN readPC[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.650 846.590 821.930 850.590 ;
    END
  END readPC[9]
  PIN sysmem_client_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 3.440 839.870 4.040 ;
    END
  END sysmem_client_ack_i
  PIN sysmem_client_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 46.960 839.870 47.560 ;
    END
  END sysmem_client_adr_o[0]
  PIN sysmem_client_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 293.800 839.870 294.400 ;
    END
  END sysmem_client_adr_o[10]
  PIN sysmem_client_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 315.560 839.870 316.160 ;
    END
  END sysmem_client_adr_o[11]
  PIN sysmem_client_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 337.320 839.870 337.920 ;
    END
  END sysmem_client_adr_o[12]
  PIN sysmem_client_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 359.080 839.870 359.680 ;
    END
  END sysmem_client_adr_o[13]
  PIN sysmem_client_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 381.520 839.870 382.120 ;
    END
  END sysmem_client_adr_o[14]
  PIN sysmem_client_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 403.280 839.870 403.880 ;
    END
  END sysmem_client_adr_o[15]
  PIN sysmem_client_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 425.040 839.870 425.640 ;
    END
  END sysmem_client_adr_o[16]
  PIN sysmem_client_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 446.800 839.870 447.400 ;
    END
  END sysmem_client_adr_o[17]
  PIN sysmem_client_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 468.560 839.870 469.160 ;
    END
  END sysmem_client_adr_o[18]
  PIN sysmem_client_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 490.320 839.870 490.920 ;
    END
  END sysmem_client_adr_o[19]
  PIN sysmem_client_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 75.520 839.870 76.120 ;
    END
  END sysmem_client_adr_o[1]
  PIN sysmem_client_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 512.080 839.870 512.680 ;
    END
  END sysmem_client_adr_o[20]
  PIN sysmem_client_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 533.840 839.870 534.440 ;
    END
  END sysmem_client_adr_o[21]
  PIN sysmem_client_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 555.600 839.870 556.200 ;
    END
  END sysmem_client_adr_o[22]
  PIN sysmem_client_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 577.360 839.870 577.960 ;
    END
  END sysmem_client_adr_o[23]
  PIN sysmem_client_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 599.120 839.870 599.720 ;
    END
  END sysmem_client_adr_o[24]
  PIN sysmem_client_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 620.880 839.870 621.480 ;
    END
  END sysmem_client_adr_o[25]
  PIN sysmem_client_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 642.640 839.870 643.240 ;
    END
  END sysmem_client_adr_o[26]
  PIN sysmem_client_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 665.080 839.870 665.680 ;
    END
  END sysmem_client_adr_o[27]
  PIN sysmem_client_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 686.840 839.870 687.440 ;
    END
  END sysmem_client_adr_o[28]
  PIN sysmem_client_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 708.600 839.870 709.200 ;
    END
  END sysmem_client_adr_o[29]
  PIN sysmem_client_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 104.760 839.870 105.360 ;
    END
  END sysmem_client_adr_o[2]
  PIN sysmem_client_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 730.360 839.870 730.960 ;
    END
  END sysmem_client_adr_o[30]
  PIN sysmem_client_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 752.120 839.870 752.720 ;
    END
  END sysmem_client_adr_o[31]
  PIN sysmem_client_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 134.000 839.870 134.600 ;
    END
  END sysmem_client_adr_o[3]
  PIN sysmem_client_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 163.240 839.870 163.840 ;
    END
  END sysmem_client_adr_o[4]
  PIN sysmem_client_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 185.000 839.870 185.600 ;
    END
  END sysmem_client_adr_o[5]
  PIN sysmem_client_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 206.760 839.870 207.360 ;
    END
  END sysmem_client_adr_o[6]
  PIN sysmem_client_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 228.520 839.870 229.120 ;
    END
  END sysmem_client_adr_o[7]
  PIN sysmem_client_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 250.280 839.870 250.880 ;
    END
  END sysmem_client_adr_o[8]
  PIN sysmem_client_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 272.040 839.870 272.640 ;
    END
  END sysmem_client_adr_o[9]
  PIN sysmem_client_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 10.240 839.870 10.840 ;
    END
  END sysmem_client_cyc_o
  PIN sysmem_client_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 53.760 839.870 54.360 ;
    END
  END sysmem_client_dat_i[0]
  PIN sysmem_client_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 301.280 839.870 301.880 ;
    END
  END sysmem_client_dat_i[10]
  PIN sysmem_client_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 323.040 839.870 323.640 ;
    END
  END sysmem_client_dat_i[11]
  PIN sysmem_client_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 344.800 839.870 345.400 ;
    END
  END sysmem_client_dat_i[12]
  PIN sysmem_client_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 366.560 839.870 367.160 ;
    END
  END sysmem_client_dat_i[13]
  PIN sysmem_client_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 388.320 839.870 388.920 ;
    END
  END sysmem_client_dat_i[14]
  PIN sysmem_client_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 410.080 839.870 410.680 ;
    END
  END sysmem_client_dat_i[15]
  PIN sysmem_client_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 431.840 839.870 432.440 ;
    END
  END sysmem_client_dat_i[16]
  PIN sysmem_client_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 453.600 839.870 454.200 ;
    END
  END sysmem_client_dat_i[17]
  PIN sysmem_client_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 476.040 839.870 476.640 ;
    END
  END sysmem_client_dat_i[18]
  PIN sysmem_client_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 497.800 839.870 498.400 ;
    END
  END sysmem_client_dat_i[19]
  PIN sysmem_client_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 83.000 839.870 83.600 ;
    END
  END sysmem_client_dat_i[1]
  PIN sysmem_client_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 519.560 839.870 520.160 ;
    END
  END sysmem_client_dat_i[20]
  PIN sysmem_client_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 541.320 839.870 541.920 ;
    END
  END sysmem_client_dat_i[21]
  PIN sysmem_client_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 563.080 839.870 563.680 ;
    END
  END sysmem_client_dat_i[22]
  PIN sysmem_client_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 584.840 839.870 585.440 ;
    END
  END sysmem_client_dat_i[23]
  PIN sysmem_client_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 606.600 839.870 607.200 ;
    END
  END sysmem_client_dat_i[24]
  PIN sysmem_client_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 628.360 839.870 628.960 ;
    END
  END sysmem_client_dat_i[25]
  PIN sysmem_client_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 650.120 839.870 650.720 ;
    END
  END sysmem_client_dat_i[26]
  PIN sysmem_client_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 671.880 839.870 672.480 ;
    END
  END sysmem_client_dat_i[27]
  PIN sysmem_client_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 693.640 839.870 694.240 ;
    END
  END sysmem_client_dat_i[28]
  PIN sysmem_client_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 715.400 839.870 716.000 ;
    END
  END sysmem_client_dat_i[29]
  PIN sysmem_client_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 112.240 839.870 112.840 ;
    END
  END sysmem_client_dat_i[2]
  PIN sysmem_client_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 737.160 839.870 737.760 ;
    END
  END sysmem_client_dat_i[30]
  PIN sysmem_client_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 759.600 839.870 760.200 ;
    END
  END sysmem_client_dat_i[31]
  PIN sysmem_client_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 141.480 839.870 142.080 ;
    END
  END sysmem_client_dat_i[3]
  PIN sysmem_client_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 170.040 839.870 170.640 ;
    END
  END sysmem_client_dat_i[4]
  PIN sysmem_client_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 192.480 839.870 193.080 ;
    END
  END sysmem_client_dat_i[5]
  PIN sysmem_client_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 214.240 839.870 214.840 ;
    END
  END sysmem_client_dat_i[6]
  PIN sysmem_client_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 236.000 839.870 236.600 ;
    END
  END sysmem_client_dat_i[7]
  PIN sysmem_client_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 257.760 839.870 258.360 ;
    END
  END sysmem_client_dat_i[8]
  PIN sysmem_client_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 279.520 839.870 280.120 ;
    END
  END sysmem_client_dat_i[9]
  PIN sysmem_client_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 61.240 839.870 61.840 ;
    END
  END sysmem_client_dat_o[0]
  PIN sysmem_client_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 308.760 839.870 309.360 ;
    END
  END sysmem_client_dat_o[10]
  PIN sysmem_client_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 330.520 839.870 331.120 ;
    END
  END sysmem_client_dat_o[11]
  PIN sysmem_client_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 352.280 839.870 352.880 ;
    END
  END sysmem_client_dat_o[12]
  PIN sysmem_client_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 374.040 839.870 374.640 ;
    END
  END sysmem_client_dat_o[13]
  PIN sysmem_client_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 395.800 839.870 396.400 ;
    END
  END sysmem_client_dat_o[14]
  PIN sysmem_client_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 417.560 839.870 418.160 ;
    END
  END sysmem_client_dat_o[15]
  PIN sysmem_client_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 439.320 839.870 439.920 ;
    END
  END sysmem_client_dat_o[16]
  PIN sysmem_client_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 461.080 839.870 461.680 ;
    END
  END sysmem_client_dat_o[17]
  PIN sysmem_client_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 482.840 839.870 483.440 ;
    END
  END sysmem_client_dat_o[18]
  PIN sysmem_client_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 504.600 839.870 505.200 ;
    END
  END sysmem_client_dat_o[19]
  PIN sysmem_client_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 90.480 839.870 91.080 ;
    END
  END sysmem_client_dat_o[1]
  PIN sysmem_client_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 526.360 839.870 526.960 ;
    END
  END sysmem_client_dat_o[20]
  PIN sysmem_client_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 548.120 839.870 548.720 ;
    END
  END sysmem_client_dat_o[21]
  PIN sysmem_client_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 570.560 839.870 571.160 ;
    END
  END sysmem_client_dat_o[22]
  PIN sysmem_client_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 592.320 839.870 592.920 ;
    END
  END sysmem_client_dat_o[23]
  PIN sysmem_client_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 614.080 839.870 614.680 ;
    END
  END sysmem_client_dat_o[24]
  PIN sysmem_client_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 635.840 839.870 636.440 ;
    END
  END sysmem_client_dat_o[25]
  PIN sysmem_client_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 657.600 839.870 658.200 ;
    END
  END sysmem_client_dat_o[26]
  PIN sysmem_client_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 679.360 839.870 679.960 ;
    END
  END sysmem_client_dat_o[27]
  PIN sysmem_client_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 701.120 839.870 701.720 ;
    END
  END sysmem_client_dat_o[28]
  PIN sysmem_client_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 722.880 839.870 723.480 ;
    END
  END sysmem_client_dat_o[29]
  PIN sysmem_client_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 119.720 839.870 120.320 ;
    END
  END sysmem_client_dat_o[2]
  PIN sysmem_client_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 744.640 839.870 745.240 ;
    END
  END sysmem_client_dat_o[30]
  PIN sysmem_client_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 766.400 839.870 767.000 ;
    END
  END sysmem_client_dat_o[31]
  PIN sysmem_client_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 148.280 839.870 148.880 ;
    END
  END sysmem_client_dat_o[3]
  PIN sysmem_client_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 177.520 839.870 178.120 ;
    END
  END sysmem_client_dat_o[4]
  PIN sysmem_client_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 199.280 839.870 199.880 ;
    END
  END sysmem_client_dat_o[5]
  PIN sysmem_client_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 221.040 839.870 221.640 ;
    END
  END sysmem_client_dat_o[6]
  PIN sysmem_client_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 242.800 839.870 243.400 ;
    END
  END sysmem_client_dat_o[7]
  PIN sysmem_client_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 264.560 839.870 265.160 ;
    END
  END sysmem_client_dat_o[8]
  PIN sysmem_client_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 287.000 839.870 287.600 ;
    END
  END sysmem_client_dat_o[9]
  PIN sysmem_client_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 17.720 839.870 18.320 ;
    END
  END sysmem_client_err_i
  PIN sysmem_client_rty_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 25.200 839.870 25.800 ;
    END
  END sysmem_client_rty_i
  PIN sysmem_client_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 68.720 839.870 69.320 ;
    END
  END sysmem_client_sel_o[0]
  PIN sysmem_client_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 97.960 839.870 98.560 ;
    END
  END sysmem_client_sel_o[1]
  PIN sysmem_client_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 126.520 839.870 127.120 ;
    END
  END sysmem_client_sel_o[2]
  PIN sysmem_client_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 155.760 839.870 156.360 ;
    END
  END sysmem_client_sel_o[3]
  PIN sysmem_client_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 32.000 839.870 32.600 ;
    END
  END sysmem_client_stb_o
  PIN sysmem_client_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 835.870 39.480 839.870 40.080 ;
    END
  END sysmem_client_we_o
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 838.000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 838.000 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 833.980 837.845 ;
      LAYER met1 ;
        RECT 0.070 10.640 838.050 841.120 ;
      LAYER met2 ;
        RECT 0.100 846.310 1.650 847.010 ;
        RECT 2.490 846.310 5.330 847.010 ;
        RECT 6.170 846.310 9.470 847.010 ;
        RECT 10.310 846.310 13.610 847.010 ;
        RECT 14.450 846.310 17.290 847.010 ;
        RECT 18.130 846.310 21.430 847.010 ;
        RECT 22.270 846.310 25.570 847.010 ;
        RECT 26.410 846.310 29.250 847.010 ;
        RECT 30.090 846.310 33.390 847.010 ;
        RECT 34.230 846.310 37.530 847.010 ;
        RECT 38.370 846.310 41.210 847.010 ;
        RECT 42.050 846.310 45.350 847.010 ;
        RECT 46.190 846.310 49.490 847.010 ;
        RECT 50.330 846.310 53.630 847.010 ;
        RECT 54.470 846.310 57.310 847.010 ;
        RECT 58.150 846.310 61.450 847.010 ;
        RECT 62.290 846.310 65.590 847.010 ;
        RECT 66.430 846.310 69.270 847.010 ;
        RECT 70.110 846.310 73.410 847.010 ;
        RECT 74.250 846.310 77.550 847.010 ;
        RECT 78.390 846.310 81.230 847.010 ;
        RECT 82.070 846.310 85.370 847.010 ;
        RECT 86.210 846.310 89.510 847.010 ;
        RECT 90.350 846.310 93.190 847.010 ;
        RECT 94.030 846.310 97.330 847.010 ;
        RECT 98.170 846.310 101.470 847.010 ;
        RECT 102.310 846.310 105.610 847.010 ;
        RECT 106.450 846.310 109.290 847.010 ;
        RECT 110.130 846.310 113.430 847.010 ;
        RECT 114.270 846.310 117.570 847.010 ;
        RECT 118.410 846.310 121.250 847.010 ;
        RECT 122.090 846.310 125.390 847.010 ;
        RECT 126.230 846.310 129.530 847.010 ;
        RECT 130.370 846.310 133.210 847.010 ;
        RECT 134.050 846.310 137.350 847.010 ;
        RECT 138.190 846.310 141.490 847.010 ;
        RECT 142.330 846.310 145.630 847.010 ;
        RECT 146.470 846.310 149.310 847.010 ;
        RECT 150.150 846.310 153.450 847.010 ;
        RECT 154.290 846.310 157.590 847.010 ;
        RECT 158.430 846.310 161.270 847.010 ;
        RECT 162.110 846.310 165.410 847.010 ;
        RECT 166.250 846.310 169.550 847.010 ;
        RECT 170.390 846.310 173.230 847.010 ;
        RECT 174.070 846.310 177.370 847.010 ;
        RECT 178.210 846.310 181.510 847.010 ;
        RECT 182.350 846.310 185.190 847.010 ;
        RECT 186.030 846.310 189.330 847.010 ;
        RECT 190.170 846.310 193.470 847.010 ;
        RECT 194.310 846.310 197.610 847.010 ;
        RECT 198.450 846.310 201.290 847.010 ;
        RECT 202.130 846.310 205.430 847.010 ;
        RECT 206.270 846.310 209.570 847.010 ;
        RECT 210.410 846.310 213.250 847.010 ;
        RECT 214.090 846.310 217.390 847.010 ;
        RECT 218.230 846.310 221.530 847.010 ;
        RECT 222.370 846.310 225.210 847.010 ;
        RECT 226.050 846.310 229.350 847.010 ;
        RECT 230.190 846.310 233.490 847.010 ;
        RECT 234.330 846.310 237.630 847.010 ;
        RECT 238.470 846.310 241.310 847.010 ;
        RECT 242.150 846.310 245.450 847.010 ;
        RECT 246.290 846.310 249.590 847.010 ;
        RECT 250.430 846.310 253.270 847.010 ;
        RECT 254.110 846.310 257.410 847.010 ;
        RECT 258.250 846.310 261.550 847.010 ;
        RECT 262.390 846.310 265.230 847.010 ;
        RECT 266.070 846.310 269.370 847.010 ;
        RECT 270.210 846.310 273.510 847.010 ;
        RECT 274.350 846.310 277.190 847.010 ;
        RECT 278.030 846.310 281.330 847.010 ;
        RECT 282.170 846.310 285.470 847.010 ;
        RECT 286.310 846.310 289.610 847.010 ;
        RECT 290.450 846.310 293.290 847.010 ;
        RECT 294.130 846.310 297.430 847.010 ;
        RECT 298.270 846.310 301.570 847.010 ;
        RECT 302.410 846.310 305.250 847.010 ;
        RECT 306.090 846.310 309.390 847.010 ;
        RECT 310.230 846.310 313.530 847.010 ;
        RECT 314.370 846.310 317.210 847.010 ;
        RECT 318.050 846.310 321.350 847.010 ;
        RECT 322.190 846.310 325.490 847.010 ;
        RECT 326.330 846.310 329.630 847.010 ;
        RECT 330.470 846.310 333.310 847.010 ;
        RECT 334.150 846.310 337.450 847.010 ;
        RECT 338.290 846.310 341.590 847.010 ;
        RECT 342.430 846.310 345.270 847.010 ;
        RECT 346.110 846.310 349.410 847.010 ;
        RECT 350.250 846.310 353.550 847.010 ;
        RECT 354.390 846.310 357.230 847.010 ;
        RECT 358.070 846.310 361.370 847.010 ;
        RECT 362.210 846.310 365.510 847.010 ;
        RECT 366.350 846.310 369.190 847.010 ;
        RECT 370.030 846.310 373.330 847.010 ;
        RECT 374.170 846.310 377.470 847.010 ;
        RECT 378.310 846.310 381.610 847.010 ;
        RECT 382.450 846.310 385.290 847.010 ;
        RECT 386.130 846.310 389.430 847.010 ;
        RECT 390.270 846.310 393.570 847.010 ;
        RECT 394.410 846.310 397.250 847.010 ;
        RECT 398.090 846.310 401.390 847.010 ;
        RECT 402.230 846.310 405.530 847.010 ;
        RECT 406.370 846.310 409.210 847.010 ;
        RECT 410.050 846.310 413.350 847.010 ;
        RECT 414.190 846.310 417.490 847.010 ;
        RECT 418.330 846.310 421.630 847.010 ;
        RECT 422.470 846.310 425.310 847.010 ;
        RECT 426.150 846.310 429.450 847.010 ;
        RECT 430.290 846.310 433.590 847.010 ;
        RECT 434.430 846.310 437.270 847.010 ;
        RECT 438.110 846.310 441.410 847.010 ;
        RECT 442.250 846.310 445.550 847.010 ;
        RECT 446.390 846.310 449.230 847.010 ;
        RECT 450.070 846.310 453.370 847.010 ;
        RECT 454.210 846.310 457.510 847.010 ;
        RECT 458.350 846.310 461.190 847.010 ;
        RECT 462.030 846.310 465.330 847.010 ;
        RECT 466.170 846.310 469.470 847.010 ;
        RECT 470.310 846.310 473.610 847.010 ;
        RECT 474.450 846.310 477.290 847.010 ;
        RECT 478.130 846.310 481.430 847.010 ;
        RECT 482.270 846.310 485.570 847.010 ;
        RECT 486.410 846.310 489.250 847.010 ;
        RECT 490.090 846.310 493.390 847.010 ;
        RECT 494.230 846.310 497.530 847.010 ;
        RECT 498.370 846.310 501.210 847.010 ;
        RECT 502.050 846.310 505.350 847.010 ;
        RECT 506.190 846.310 509.490 847.010 ;
        RECT 510.330 846.310 513.170 847.010 ;
        RECT 514.010 846.310 517.310 847.010 ;
        RECT 518.150 846.310 521.450 847.010 ;
        RECT 522.290 846.310 525.590 847.010 ;
        RECT 526.430 846.310 529.270 847.010 ;
        RECT 530.110 846.310 533.410 847.010 ;
        RECT 534.250 846.310 537.550 847.010 ;
        RECT 538.390 846.310 541.230 847.010 ;
        RECT 542.070 846.310 545.370 847.010 ;
        RECT 546.210 846.310 549.510 847.010 ;
        RECT 550.350 846.310 553.190 847.010 ;
        RECT 554.030 846.310 557.330 847.010 ;
        RECT 558.170 846.310 561.470 847.010 ;
        RECT 562.310 846.310 565.610 847.010 ;
        RECT 566.450 846.310 569.290 847.010 ;
        RECT 570.130 846.310 573.430 847.010 ;
        RECT 574.270 846.310 577.570 847.010 ;
        RECT 578.410 846.310 581.250 847.010 ;
        RECT 582.090 846.310 585.390 847.010 ;
        RECT 586.230 846.310 589.530 847.010 ;
        RECT 590.370 846.310 593.210 847.010 ;
        RECT 594.050 846.310 597.350 847.010 ;
        RECT 598.190 846.310 601.490 847.010 ;
        RECT 602.330 846.310 605.170 847.010 ;
        RECT 606.010 846.310 609.310 847.010 ;
        RECT 610.150 846.310 613.450 847.010 ;
        RECT 614.290 846.310 617.590 847.010 ;
        RECT 618.430 846.310 621.270 847.010 ;
        RECT 622.110 846.310 625.410 847.010 ;
        RECT 626.250 846.310 629.550 847.010 ;
        RECT 630.390 846.310 633.230 847.010 ;
        RECT 634.070 846.310 637.370 847.010 ;
        RECT 638.210 846.310 641.510 847.010 ;
        RECT 642.350 846.310 645.190 847.010 ;
        RECT 646.030 846.310 649.330 847.010 ;
        RECT 650.170 846.310 653.470 847.010 ;
        RECT 654.310 846.310 657.610 847.010 ;
        RECT 658.450 846.310 661.290 847.010 ;
        RECT 662.130 846.310 665.430 847.010 ;
        RECT 666.270 846.310 669.570 847.010 ;
        RECT 670.410 846.310 673.250 847.010 ;
        RECT 674.090 846.310 677.390 847.010 ;
        RECT 678.230 846.310 681.530 847.010 ;
        RECT 682.370 846.310 685.210 847.010 ;
        RECT 686.050 846.310 689.350 847.010 ;
        RECT 690.190 846.310 693.490 847.010 ;
        RECT 694.330 846.310 697.170 847.010 ;
        RECT 698.010 846.310 701.310 847.010 ;
        RECT 702.150 846.310 705.450 847.010 ;
        RECT 706.290 846.310 709.590 847.010 ;
        RECT 710.430 846.310 713.270 847.010 ;
        RECT 714.110 846.310 717.410 847.010 ;
        RECT 718.250 846.310 721.550 847.010 ;
        RECT 722.390 846.310 725.230 847.010 ;
        RECT 726.070 846.310 729.370 847.010 ;
        RECT 730.210 846.310 733.510 847.010 ;
        RECT 734.350 846.310 737.190 847.010 ;
        RECT 738.030 846.310 741.330 847.010 ;
        RECT 742.170 846.310 745.470 847.010 ;
        RECT 746.310 846.310 749.610 847.010 ;
        RECT 750.450 846.310 753.290 847.010 ;
        RECT 754.130 846.310 757.430 847.010 ;
        RECT 758.270 846.310 761.570 847.010 ;
        RECT 762.410 846.310 765.250 847.010 ;
        RECT 766.090 846.310 769.390 847.010 ;
        RECT 770.230 846.310 773.530 847.010 ;
        RECT 774.370 846.310 777.210 847.010 ;
        RECT 778.050 846.310 781.350 847.010 ;
        RECT 782.190 846.310 785.490 847.010 ;
        RECT 786.330 846.310 789.170 847.010 ;
        RECT 790.010 846.310 793.310 847.010 ;
        RECT 794.150 846.310 797.450 847.010 ;
        RECT 798.290 846.310 801.590 847.010 ;
        RECT 802.430 846.310 805.270 847.010 ;
        RECT 806.110 846.310 809.410 847.010 ;
        RECT 810.250 846.310 813.550 847.010 ;
        RECT 814.390 846.310 817.230 847.010 ;
        RECT 818.070 846.310 821.370 847.010 ;
        RECT 822.210 846.310 825.510 847.010 ;
        RECT 826.350 846.310 829.190 847.010 ;
        RECT 830.030 846.310 833.330 847.010 ;
        RECT 834.170 846.310 837.470 847.010 ;
        RECT 0.100 4.280 838.020 846.310 ;
        RECT 0.100 3.555 83.530 4.280 ;
        RECT 84.370 3.555 251.430 4.280 ;
        RECT 252.270 3.555 419.330 4.280 ;
        RECT 420.170 3.555 587.230 4.280 ;
        RECT 588.070 3.555 755.130 4.280 ;
        RECT 755.970 3.555 838.020 4.280 ;
      LAYER met3 ;
        RECT 4.000 846.240 835.470 847.090 ;
        RECT 4.000 840.160 835.870 846.240 ;
        RECT 4.000 838.760 835.470 840.160 ;
        RECT 4.000 832.680 835.870 838.760 ;
        RECT 4.000 831.280 835.470 832.680 ;
        RECT 4.000 825.880 835.870 831.280 ;
        RECT 4.000 824.480 835.470 825.880 ;
        RECT 4.000 818.400 835.870 824.480 ;
        RECT 4.400 817.000 835.470 818.400 ;
        RECT 4.000 810.920 835.870 817.000 ;
        RECT 4.000 809.520 835.470 810.920 ;
        RECT 4.000 804.120 835.870 809.520 ;
        RECT 4.000 802.720 835.470 804.120 ;
        RECT 4.000 796.640 835.870 802.720 ;
        RECT 4.000 795.240 835.470 796.640 ;
        RECT 4.000 789.160 835.870 795.240 ;
        RECT 4.000 787.760 835.470 789.160 ;
        RECT 4.000 782.360 835.870 787.760 ;
        RECT 4.000 780.960 835.470 782.360 ;
        RECT 4.000 774.880 835.870 780.960 ;
        RECT 4.000 773.480 835.470 774.880 ;
        RECT 4.000 767.400 835.870 773.480 ;
        RECT 4.000 766.000 835.470 767.400 ;
        RECT 4.000 760.600 835.870 766.000 ;
        RECT 4.000 759.200 835.470 760.600 ;
        RECT 4.000 753.120 835.870 759.200 ;
        RECT 4.400 751.720 835.470 753.120 ;
        RECT 4.000 745.640 835.870 751.720 ;
        RECT 4.000 744.240 835.470 745.640 ;
        RECT 4.000 738.160 835.870 744.240 ;
        RECT 4.000 736.760 835.470 738.160 ;
        RECT 4.000 731.360 835.870 736.760 ;
        RECT 4.000 729.960 835.470 731.360 ;
        RECT 4.000 723.880 835.870 729.960 ;
        RECT 4.000 722.480 835.470 723.880 ;
        RECT 4.000 716.400 835.870 722.480 ;
        RECT 4.000 715.000 835.470 716.400 ;
        RECT 4.000 709.600 835.870 715.000 ;
        RECT 4.000 708.200 835.470 709.600 ;
        RECT 4.000 702.120 835.870 708.200 ;
        RECT 4.000 700.720 835.470 702.120 ;
        RECT 4.000 694.640 835.870 700.720 ;
        RECT 4.000 693.240 835.470 694.640 ;
        RECT 4.000 687.840 835.870 693.240 ;
        RECT 4.400 686.440 835.470 687.840 ;
        RECT 4.000 680.360 835.870 686.440 ;
        RECT 4.000 678.960 835.470 680.360 ;
        RECT 4.000 672.880 835.870 678.960 ;
        RECT 4.000 671.480 835.470 672.880 ;
        RECT 4.000 666.080 835.870 671.480 ;
        RECT 4.000 664.680 835.470 666.080 ;
        RECT 4.000 658.600 835.870 664.680 ;
        RECT 4.000 657.200 835.470 658.600 ;
        RECT 4.000 651.120 835.870 657.200 ;
        RECT 4.000 649.720 835.470 651.120 ;
        RECT 4.000 643.640 835.870 649.720 ;
        RECT 4.000 642.240 835.470 643.640 ;
        RECT 4.000 636.840 835.870 642.240 ;
        RECT 4.000 635.440 835.470 636.840 ;
        RECT 4.000 629.360 835.870 635.440 ;
        RECT 4.000 627.960 835.470 629.360 ;
        RECT 4.000 622.560 835.870 627.960 ;
        RECT 4.400 621.880 835.870 622.560 ;
        RECT 4.400 621.160 835.470 621.880 ;
        RECT 4.000 620.480 835.470 621.160 ;
        RECT 4.000 615.080 835.870 620.480 ;
        RECT 4.000 613.680 835.470 615.080 ;
        RECT 4.000 607.600 835.870 613.680 ;
        RECT 4.000 606.200 835.470 607.600 ;
        RECT 4.000 600.120 835.870 606.200 ;
        RECT 4.000 598.720 835.470 600.120 ;
        RECT 4.000 593.320 835.870 598.720 ;
        RECT 4.000 591.920 835.470 593.320 ;
        RECT 4.000 585.840 835.870 591.920 ;
        RECT 4.000 584.440 835.470 585.840 ;
        RECT 4.000 578.360 835.870 584.440 ;
        RECT 4.000 576.960 835.470 578.360 ;
        RECT 4.000 571.560 835.870 576.960 ;
        RECT 4.000 570.160 835.470 571.560 ;
        RECT 4.000 564.080 835.870 570.160 ;
        RECT 4.000 562.680 835.470 564.080 ;
        RECT 4.000 556.600 835.870 562.680 ;
        RECT 4.400 555.200 835.470 556.600 ;
        RECT 4.000 549.120 835.870 555.200 ;
        RECT 4.000 547.720 835.470 549.120 ;
        RECT 4.000 542.320 835.870 547.720 ;
        RECT 4.000 540.920 835.470 542.320 ;
        RECT 4.000 534.840 835.870 540.920 ;
        RECT 4.000 533.440 835.470 534.840 ;
        RECT 4.000 527.360 835.870 533.440 ;
        RECT 4.000 525.960 835.470 527.360 ;
        RECT 4.000 520.560 835.870 525.960 ;
        RECT 4.000 519.160 835.470 520.560 ;
        RECT 4.000 513.080 835.870 519.160 ;
        RECT 4.000 511.680 835.470 513.080 ;
        RECT 4.000 505.600 835.870 511.680 ;
        RECT 4.000 504.200 835.470 505.600 ;
        RECT 4.000 498.800 835.870 504.200 ;
        RECT 4.000 497.400 835.470 498.800 ;
        RECT 4.000 491.320 835.870 497.400 ;
        RECT 4.400 489.920 835.470 491.320 ;
        RECT 4.000 483.840 835.870 489.920 ;
        RECT 4.000 482.440 835.470 483.840 ;
        RECT 4.000 477.040 835.870 482.440 ;
        RECT 4.000 475.640 835.470 477.040 ;
        RECT 4.000 469.560 835.870 475.640 ;
        RECT 4.000 468.160 835.470 469.560 ;
        RECT 4.000 462.080 835.870 468.160 ;
        RECT 4.000 460.680 835.470 462.080 ;
        RECT 4.000 454.600 835.870 460.680 ;
        RECT 4.000 453.200 835.470 454.600 ;
        RECT 4.000 447.800 835.870 453.200 ;
        RECT 4.000 446.400 835.470 447.800 ;
        RECT 4.000 440.320 835.870 446.400 ;
        RECT 4.000 438.920 835.470 440.320 ;
        RECT 4.000 432.840 835.870 438.920 ;
        RECT 4.000 431.440 835.470 432.840 ;
        RECT 4.000 426.040 835.870 431.440 ;
        RECT 4.400 424.640 835.470 426.040 ;
        RECT 4.000 418.560 835.870 424.640 ;
        RECT 4.000 417.160 835.470 418.560 ;
        RECT 4.000 411.080 835.870 417.160 ;
        RECT 4.000 409.680 835.470 411.080 ;
        RECT 4.000 404.280 835.870 409.680 ;
        RECT 4.000 402.880 835.470 404.280 ;
        RECT 4.000 396.800 835.870 402.880 ;
        RECT 4.000 395.400 835.470 396.800 ;
        RECT 4.000 389.320 835.870 395.400 ;
        RECT 4.000 387.920 835.470 389.320 ;
        RECT 4.000 382.520 835.870 387.920 ;
        RECT 4.000 381.120 835.470 382.520 ;
        RECT 4.000 375.040 835.870 381.120 ;
        RECT 4.000 373.640 835.470 375.040 ;
        RECT 4.000 367.560 835.870 373.640 ;
        RECT 4.000 366.160 835.470 367.560 ;
        RECT 4.000 360.760 835.870 366.160 ;
        RECT 4.400 360.080 835.870 360.760 ;
        RECT 4.400 359.360 835.470 360.080 ;
        RECT 4.000 358.680 835.470 359.360 ;
        RECT 4.000 353.280 835.870 358.680 ;
        RECT 4.000 351.880 835.470 353.280 ;
        RECT 4.000 345.800 835.870 351.880 ;
        RECT 4.000 344.400 835.470 345.800 ;
        RECT 4.000 338.320 835.870 344.400 ;
        RECT 4.000 336.920 835.470 338.320 ;
        RECT 4.000 331.520 835.870 336.920 ;
        RECT 4.000 330.120 835.470 331.520 ;
        RECT 4.000 324.040 835.870 330.120 ;
        RECT 4.000 322.640 835.470 324.040 ;
        RECT 4.000 316.560 835.870 322.640 ;
        RECT 4.000 315.160 835.470 316.560 ;
        RECT 4.000 309.760 835.870 315.160 ;
        RECT 4.000 308.360 835.470 309.760 ;
        RECT 4.000 302.280 835.870 308.360 ;
        RECT 4.000 300.880 835.470 302.280 ;
        RECT 4.000 294.800 835.870 300.880 ;
        RECT 4.400 293.400 835.470 294.800 ;
        RECT 4.000 288.000 835.870 293.400 ;
        RECT 4.000 286.600 835.470 288.000 ;
        RECT 4.000 280.520 835.870 286.600 ;
        RECT 4.000 279.120 835.470 280.520 ;
        RECT 4.000 273.040 835.870 279.120 ;
        RECT 4.000 271.640 835.470 273.040 ;
        RECT 4.000 265.560 835.870 271.640 ;
        RECT 4.000 264.160 835.470 265.560 ;
        RECT 4.000 258.760 835.870 264.160 ;
        RECT 4.000 257.360 835.470 258.760 ;
        RECT 4.000 251.280 835.870 257.360 ;
        RECT 4.000 249.880 835.470 251.280 ;
        RECT 4.000 243.800 835.870 249.880 ;
        RECT 4.000 242.400 835.470 243.800 ;
        RECT 4.000 237.000 835.870 242.400 ;
        RECT 4.000 235.600 835.470 237.000 ;
        RECT 4.000 229.520 835.870 235.600 ;
        RECT 4.400 228.120 835.470 229.520 ;
        RECT 4.000 222.040 835.870 228.120 ;
        RECT 4.000 220.640 835.470 222.040 ;
        RECT 4.000 215.240 835.870 220.640 ;
        RECT 4.000 213.840 835.470 215.240 ;
        RECT 4.000 207.760 835.870 213.840 ;
        RECT 4.000 206.360 835.470 207.760 ;
        RECT 4.000 200.280 835.870 206.360 ;
        RECT 4.000 198.880 835.470 200.280 ;
        RECT 4.000 193.480 835.870 198.880 ;
        RECT 4.000 192.080 835.470 193.480 ;
        RECT 4.000 186.000 835.870 192.080 ;
        RECT 4.000 184.600 835.470 186.000 ;
        RECT 4.000 178.520 835.870 184.600 ;
        RECT 4.000 177.120 835.470 178.520 ;
        RECT 4.000 171.040 835.870 177.120 ;
        RECT 4.000 169.640 835.470 171.040 ;
        RECT 4.000 164.240 835.870 169.640 ;
        RECT 4.400 162.840 835.470 164.240 ;
        RECT 4.000 156.760 835.870 162.840 ;
        RECT 4.000 155.360 835.470 156.760 ;
        RECT 4.000 149.280 835.870 155.360 ;
        RECT 4.000 147.880 835.470 149.280 ;
        RECT 4.000 142.480 835.870 147.880 ;
        RECT 4.000 141.080 835.470 142.480 ;
        RECT 4.000 135.000 835.870 141.080 ;
        RECT 4.000 133.600 835.470 135.000 ;
        RECT 4.000 127.520 835.870 133.600 ;
        RECT 4.000 126.120 835.470 127.520 ;
        RECT 4.000 120.720 835.870 126.120 ;
        RECT 4.000 119.320 835.470 120.720 ;
        RECT 4.000 113.240 835.870 119.320 ;
        RECT 4.000 111.840 835.470 113.240 ;
        RECT 4.000 105.760 835.870 111.840 ;
        RECT 4.000 104.360 835.470 105.760 ;
        RECT 4.000 98.960 835.870 104.360 ;
        RECT 4.400 97.560 835.470 98.960 ;
        RECT 4.000 91.480 835.870 97.560 ;
        RECT 4.000 90.080 835.470 91.480 ;
        RECT 4.000 84.000 835.870 90.080 ;
        RECT 4.000 82.600 835.470 84.000 ;
        RECT 4.000 76.520 835.870 82.600 ;
        RECT 4.000 75.120 835.470 76.520 ;
        RECT 4.000 69.720 835.870 75.120 ;
        RECT 4.000 68.320 835.470 69.720 ;
        RECT 4.000 62.240 835.870 68.320 ;
        RECT 4.000 60.840 835.470 62.240 ;
        RECT 4.000 54.760 835.870 60.840 ;
        RECT 4.000 53.360 835.470 54.760 ;
        RECT 4.000 47.960 835.870 53.360 ;
        RECT 4.000 46.560 835.470 47.960 ;
        RECT 4.000 40.480 835.870 46.560 ;
        RECT 4.000 39.080 835.470 40.480 ;
        RECT 4.000 33.680 835.870 39.080 ;
        RECT 4.400 33.000 835.870 33.680 ;
        RECT 4.400 32.280 835.470 33.000 ;
        RECT 4.000 31.600 835.470 32.280 ;
        RECT 4.000 26.200 835.870 31.600 ;
        RECT 4.000 24.800 835.470 26.200 ;
        RECT 4.000 18.720 835.870 24.800 ;
        RECT 4.000 17.320 835.470 18.720 ;
        RECT 4.000 11.240 835.870 17.320 ;
        RECT 4.000 9.840 835.470 11.240 ;
        RECT 4.000 4.440 835.870 9.840 ;
        RECT 4.000 3.575 835.470 4.440 ;
      LAYER met4 ;
        RECT 96.895 18.535 97.440 822.625 ;
        RECT 99.840 18.535 174.240 822.625 ;
        RECT 176.640 18.535 251.040 822.625 ;
        RECT 253.440 18.535 327.840 822.625 ;
        RECT 330.240 18.535 404.640 822.625 ;
        RECT 407.040 18.535 481.440 822.625 ;
        RECT 483.840 18.535 558.240 822.625 ;
        RECT 560.640 18.535 635.040 822.625 ;
        RECT 637.440 18.535 711.840 822.625 ;
        RECT 714.240 18.535 788.640 822.625 ;
        RECT 791.040 18.535 828.625 822.625 ;
  END
END mkLanaiCPU
END LIBRARY

